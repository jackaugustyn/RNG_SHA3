`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/28/2023 02:35:20 PM
// Design Name: 
// Module Name: AdaptiveProportionTest
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module AdaptiveProportionTest(
    input wire[1023:0] random_bits,
    input wire[9:0] index_of_last_bit,
    output wire failure
    );
    
    assign failure = (
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-0)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-2)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-3)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-4)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-5)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-6)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-7)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-8)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-9)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-10)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-11)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-12)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-13)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-14)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-15)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-16)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-17)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-18)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-19)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-20)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-21)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-22)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-23)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-24)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-25)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-26)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-27)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-28)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-29)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-30)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-31)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-32)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-33)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-34)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-35)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-36)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-37)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-38)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-39)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-40)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-41)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-42)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-43)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-44)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-45)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-46)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-47)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-48)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-49)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-50)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-51)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-52)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-53)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-54)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-55)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-56)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-57)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-58)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-59)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-60)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-61)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-62)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-63)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-64)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-65)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-66)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-67)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-68)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-69)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-70)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-71)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-72)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-73)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-74)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-75)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-76)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-77)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-78)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-79)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-80)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-81)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-82)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-83)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-84)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-85)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-86)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-87)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-88)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-89)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-90)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-91)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-92)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-93)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-94)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-95)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-96)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-97)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-98)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-99)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-100)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-101)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-102)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-103)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-104)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-105)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-106)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-107)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-108)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-109)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-110)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-111)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-112)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-113)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-114)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-115)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-116)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-117)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-118)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-119)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-120)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-121)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-122)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-123)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-124)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-125)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-126)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-127)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-128)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-129)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-130)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-131)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-132)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-133)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-134)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-135)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-136)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-137)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-138)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-139)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-140)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-141)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-142)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-143)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-144)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-145)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-146)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-147)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-148)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-149)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-150)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-151)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-152)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-153)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-154)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-155)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-156)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-157)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-158)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-159)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-160)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-161)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-162)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-163)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-164)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-165)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-166)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-167)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-168)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-169)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-170)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-171)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-172)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-173)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-174)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-175)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-176)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-177)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-178)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-179)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-180)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-181)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-182)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-183)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-184)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-185)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-186)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-187)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-188)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-189)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-190)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-191)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-192)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-193)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-194)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-195)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-196)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-197)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-198)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-199)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-200)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-201)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-202)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-203)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-204)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-205)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-206)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-207)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-208)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-209)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-210)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-211)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-212)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-213)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-214)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-215)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-216)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-217)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-218)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-219)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-220)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-221)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-222)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-223)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-224)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-225)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-226)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-227)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-228)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-229)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-230)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-231)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-232)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-233)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-234)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-235)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-236)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-237)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-238)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-239)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-240)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-241)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-242)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-243)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-244)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-245)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-246)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-247)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-248)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-249)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-250)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-251)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-252)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-253)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-254)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-255)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-256)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-257)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-258)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-259)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-260)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-261)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-262)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-263)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-264)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-265)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-266)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-267)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-268)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-269)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-270)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-271)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-272)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-273)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-274)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-275)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-276)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-277)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-278)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-279)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-280)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-281)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-282)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-283)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-284)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-285)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-286)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-287)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-288)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-289)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-290)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-291)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-292)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-293)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-294)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-295)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-296)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-297)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-298)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-299)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-300)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-301)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-302)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-303)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-304)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-305)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-306)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-307)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-308)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-309)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-310)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-311)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-312)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-313)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-314)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-315)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-316)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-317)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-318)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-319)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-320)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-321)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-322)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-323)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-324)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-325)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-326)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-327)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-328)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-329)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-330)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-331)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-332)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-333)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-334)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-335)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-336)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-337)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-338)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-339)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-340)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-341)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-342)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-343)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-344)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-345)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-346)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-347)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-348)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-349)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-350)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-351)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-352)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-353)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-354)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-355)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-356)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-357)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-358)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-359)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-360)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-361)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-362)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-363)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-364)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-365)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-366)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-367)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-368)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-369)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-370)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-371)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-372)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-373)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-374)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-375)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-376)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-377)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-378)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-379)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-380)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-381)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-382)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-383)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-384)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-385)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-386)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-387)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-388)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-389)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-390)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-391)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-392)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-393)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-394)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-395)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-396)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-397)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-398)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-399)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-400)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-401)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-402)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-403)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-404)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-405)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-406)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-407)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-408)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-409)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-410)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-411)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-412)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-413)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-414)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-415)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-416)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-417)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-418)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-419)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-420)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-421)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-422)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-423)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-424)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-425)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-426)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-427)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-428)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-429)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-430)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-431)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-432)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-433)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-434)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-435)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-436)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-437)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-438)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-439)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-440)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-441)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-442)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-443)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-444)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-445)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-446)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-447)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-448)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-449)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-450)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-451)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-452)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-453)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-454)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-455)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-456)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-457)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-458)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-459)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-460)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-461)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-462)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-463)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-464)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-465)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-466)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-467)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-468)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-469)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-470)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-471)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-472)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-473)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-474)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-475)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-476)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-477)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-478)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-479)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-480)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-481)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-482)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-483)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-484)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-485)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-486)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-487)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-488)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-489)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-490)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-491)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-492)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-493)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-494)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-495)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-496)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-497)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-498)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-499)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-500)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-501)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-502)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-503)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-504)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-505)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-506)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-507)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-508)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-509)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-510)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-511)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-512)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-513)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-514)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-515)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-516)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-517)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-518)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-519)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-520)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-521)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-522)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-523)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-524)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-525)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-526)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-527)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-528)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-529)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-530)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-531)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-532)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-533)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-534)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-535)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-536)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-537)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-538)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-539)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-540)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-541)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-542)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-543)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-544)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-545)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-546)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-547)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-548)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-549)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-550)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-551)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-552)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-553)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-554)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-555)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-556)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-557)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-558)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-559)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-560)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-561)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-562)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-563)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-564)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-565)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-566)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-567)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-568)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-569)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-570)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-571)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-572)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-573)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-574)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-575)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-576)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-577)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-578)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-579)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-580)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-581)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-582)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-583)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-584)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-585)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-586)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-587)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-588)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-589)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-590)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-591)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-592)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-593)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-594)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-595)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-596)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-597)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-598)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-599)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-600)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-601)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-602)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-603)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-604)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-605)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-606)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-607)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-608)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-609)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-610)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-611)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-612)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-613)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-614)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-615)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-616)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-617)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-618)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-619)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-620)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-621)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-622)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-623)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-624)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-625)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-626)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-627)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-628)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-629)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-630)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-631)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-632)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-633)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-634)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-635)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-636)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-637)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-638)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-639)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-640)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-641)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-642)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-643)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-644)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-645)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-646)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-647)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-648)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-649)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-650)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-651)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-652)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-653)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-654)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-655)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-656)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-657)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-658)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-659)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-660)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-661)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-662)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-663)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-664)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-665)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-666)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-667)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-668)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-669)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-670)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-671)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-672)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-673)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-674)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-675)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-676)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-677)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-678)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-679)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-680)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-681)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-682)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-683)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-684)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-685)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-686)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-687)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-688)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-689)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-690)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-691)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-692)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-693)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-694)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-695)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-696)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-697)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-698)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-699)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-700)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-701)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-702)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-703)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-704)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-705)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-706)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-707)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-708)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-709)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-710)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-711)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-712)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-713)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-714)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-715)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-716)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-717)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-718)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-719)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-720)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-721)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-722)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-723)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-724)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-725)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-726)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-727)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-728)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-729)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-730)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-731)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-732)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-733)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-734)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-735)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-736)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-737)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-738)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-739)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-740)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-741)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-742)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-743)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-744)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-745)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-746)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-747)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-748)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-749)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-750)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-751)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-752)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-753)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-754)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-755)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-756)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-757)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-758)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-759)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-760)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-761)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-762)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-763)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-764)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-765)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-766)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-767)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-768)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-769)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-770)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-771)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-772)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-773)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-774)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-775)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-776)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-777)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-778)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-779)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-780)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-781)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-782)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-783)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-784)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-785)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-786)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-787)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-788)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-789)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-790)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-791)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-792)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-793)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-794)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-795)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-796)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-797)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-798)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-799)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-800)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-801)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-802)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-803)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-804)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-805)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-806)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-807)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-808)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-809)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-810)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-811)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-812)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-813)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-814)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-815)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-816)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-817)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-818)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-819)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-820)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-821)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-822)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-823)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-824)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-825)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-826)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-827)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-828)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-829)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-830)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-831)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-832)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-833)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-834)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-835)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-836)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-837)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-838)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-839)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-840)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-841)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-842)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-843)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-844)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-845)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-846)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-847)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-848)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-849)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-850)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-851)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-852)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-853)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-854)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-855)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-856)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-857)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-858)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-859)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-860)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-861)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-862)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-863)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-864)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-865)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-866)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-867)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-868)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-869)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-870)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-871)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-872)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-873)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-874)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-875)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-876)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-877)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-878)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-879)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-880)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-881)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-882)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-883)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-884)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-885)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-886)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-887)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-888)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-889)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-890)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-891)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-892)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-893)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-894)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-895)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-896)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-897)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-898)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-899)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-900)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-901)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-902)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-903)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-904)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-905)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-906)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-907)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-908)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-909)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-910)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-911)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-912)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-913)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-914)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-915)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-916)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-917)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-918)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-919)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-920)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-921)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-922)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-923)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-924)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-925)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-926)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-927)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-928)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-929)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-930)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-931)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-932)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-933)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-934)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-935)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-936)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-937)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-938)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-939)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-940)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-941)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-942)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-943)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-944)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-945)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-946)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-947)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-948)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-949)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-950)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-951)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-952)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-953)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-954)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-955)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-956)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-957)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-958)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-959)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-960)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-961)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-962)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-963)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-964)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-965)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-966)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-967)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-968)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-969)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-970)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-971)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-972)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-973)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-974)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-975)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-976)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-977)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-978)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-979)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-980)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-981)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-982)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-983)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-984)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-985)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-986)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-987)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-988)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-989)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-990)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-991)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-992)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-993)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-994)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-995)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-996)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-997)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-998)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-999)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1000)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1001)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1002)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1003)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1004)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1005)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1006)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1007)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1008)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1009)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1010)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1011)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1012)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1013)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1014)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1015)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1016)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1017)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1018)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1019)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1020)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1021)% 1024]) +
        (random_bits[(index_of_last_bit - 1023) % 1024] == random_bits[(index_of_last_bit-1022)% 1024])
    ) > 589 ? 1 : 0; 

    
endmodule
