`default_nettype wire
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/27/2023 01:46:18 PM
// Design Name: 
// Module Name: FiGaRO_SHA3
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module FiGaRO_SHA3(
    input  wire reset,
    input  wire enable,
    input  wire clk,
    output reg ready,
    input  wire[10:0] ADDR,
    output reg[31:0] DATA_OUT
    );
    
  parameter CHUNK_SIZE = 1023;//32767;
  parameter NUMBER_OF_WORDS_SHA3INIT = CHUNK_SIZE / 32;
    
  parameter ADDR_CTRLADDR_CTRL        = 8'h08;
  parameter CTRL_INIT_VALUE  = 8'h01;
  parameter CTRL_NEXT_VALUE  = 8'h02;
  parameter CTRL_MODE_VALUE  = 8'h04;
  
  parameter ADDR_BLOCK0    = 6'h00;
  parameter ADDR_BLOCK1    = 6'h01;
  parameter ADDR_BLOCK2    = 6'h02;
  parameter ADDR_BLOCK3    = 6'h03;
  parameter ADDR_BLOCK4    = 6'h04;
  parameter ADDR_BLOCK5    = 6'h05;
  parameter ADDR_BLOCK6    = 6'h06;
  parameter ADDR_BLOCK7    = 6'h07;
  parameter ADDR_BLOCK8    = 6'h08;
  parameter ADDR_BLOCK9    = 6'h09;
  parameter ADDR_BLOCK10   = 6'h0a;
  parameter ADDR_BLOCK11   = 6'h0b;
  parameter ADDR_BLOCK12   = 6'h0c;
  parameter ADDR_BLOCK13   = 6'h0d;
  parameter ADDR_BLOCK14   = 6'h0e;
  parameter ADDR_BLOCK15   = 6'h0f;
  parameter ADDR_BLOCK16   = 6'h10;
  parameter ADDR_BLOCK17   = 6'h11;
  parameter ADDR_BLOCK18   = 6'h12;
  parameter ADDR_BLOCK19   = 6'h13;
  parameter ADDR_BLOCK20   = 6'h14;
  parameter ADDR_BLOCK21   = 6'h15;
  parameter ADDR_BLOCK22   = 6'h16;
  parameter ADDR_BLOCK23   = 6'h17;
  parameter ADDR_BLOCK24   = 6'h18;
  parameter ADDR_BLOCK25   = 6'h19;
  parameter ADDR_BLOCK26   = 6'h1a;
  parameter ADDR_BLOCK27   = 6'h1b;
  parameter ADDR_BLOCK28   = 6'h1c;
  parameter ADDR_BLOCK29   = 6'h1d;
  parameter ADDR_BLOCK30   = 6'h1e;
  parameter ADDR_BLOCK31   = 6'h1f;
  parameter ADDR_BLOCK32   = 6'h20;
  parameter ADDR_BLOCK33   = 6'h21;
  parameter ADDR_BLOCK34   = 6'h22;
  parameter ADDR_BLOCK35   = 6'h23;
  parameter ADDR_BLOCK36   = 6'h24;
  parameter ADDR_BLOCK37   = 6'h25;
  parameter ADDR_BLOCK38   = 6'h26;
  parameter ADDR_BLOCK39   = 6'h27;
  parameter ADDR_BLOCK40   = 6'h28;
  parameter ADDR_BLOCK41   = 6'h29;
  parameter ADDR_BLOCK42   = 6'h2a;
  parameter ADDR_BLOCK43   = 6'h2b;
  parameter ADDR_BLOCK44   = 6'h2c;
  parameter ADDR_BLOCK45   = 6'h2d;
  parameter ADDR_BLOCK46   = 6'h2e;
  parameter ADDR_BLOCK47   = 6'h2f;
  parameter ADDR_BLOCK48   = 6'h30;
  parameter ADDR_BLOCK49   = 6'h31;
  parameter ADDR_BLOCK50   = 6'h32;

  parameter ADDR_DIGEST0   = 6'h40;
  parameter ADDR_DIGEST1   = 6'h41;
  parameter ADDR_DIGEST2   = 6'h42;
  parameter ADDR_DIGEST3   = 6'h43;
  parameter ADDR_DIGEST4   = 6'h44;
  parameter ADDR_DIGEST5   = 6'h45;
  parameter ADDR_DIGEST6   = 6'h46;
  parameter ADDR_DIGEST7   = 6'h47;
  parameter ADDR_DIGEST8   = 6'h48;
  parameter ADDR_DIGEST9   = 6'h49;
  parameter ADDR_DIGESTA   = 6'h4a;
  parameter ADDR_DIGESTB   = 6'h4b;
  parameter ADDR_DIGESTC   = 6'h4c;
  parameter ADDR_DIGESTD   = 6'h4d;
  parameter ADDR_DIGESTE   = 6'h4e;
  parameter ADDR_DIGESTF   = 6'h4f;

    
localparam [3:0]
    starting                = 4'b0000,
    generating              = 4'b0001,
    generated               = 4'b0010,
    writing_to_sha          = 4'b0011,
    writed_to_sha           = 4'b0100,
    generating_hash         = 4'b0101,
    hash_generated          = 4'b0110,
    final_hash_generation   = 4'b0111,
    final_hash_generated    = 4'b1000,
    saving_hash             = 4'b1001,
    saved_hash              = 4'b1010,
    increment_counter       = 4'b1011,
    sending_data            = 4'b1100,
    data_sended             = 4'b1101;


    
reg[3:0] state;

//reg[33023:0] random_bits;
reg[1023:0] random_bits;
reg[16:0] generated_bits_counter;

reg[9:0] writed_words_counter;

reg[5:0] generating_hash_counter;

wire[9:0] writed_words_counter_wire;

reg[3:0] readed_words_counter; // zlicza słowa odczytane ze skrótu

reg          sha3_init;
reg          sha3_next;
wire          sha3_ready;
reg          sha3_we;
reg[7 : 0]   sha3_address;
reg[31 : 0]  sha3_din;
wire[31 : 0]  sha3_dout;

reg [511 : 0] digest_data;


    
//RANDOM GENERATORS     
wire gen1_out, gen2_out;//, gen3_out, gen4_out, gen5_out, gen6_out, gen7_out, gen8_out;
wire random_out;
    
FiGaRO generator1(.clk(clk), .dff_en(enable), .en(enable), .random_out(gen1_out));
FiGaRO generator2(.clk(clk), .dff_en(enable), .en(enable), .random_out(gen2_out));
// FiGaRO generator3(.clk(clk), .dff_en(enable), .en(enable), .random_out(gen3_out));
// FiGaRO generator4(.clk(clk), .dff_en(enable), .en(enable), .random_out(gen4_out));
// FiGaRO generator5(.clk(clk), .dff_en(enable), .en(enable), .random_out(gen5_out));
// FiGaRO generator6(.clk(clk), .dff_en(enable), .en(enable), .random_out(gen6_out));
// FiGaRO generator7(.clk(clk), .dff_en(enable), .en(enable), .random_out(gen7_out));
// FiGaRO generator8(.clk(clk), .dff_en(enable), .en(enable), .random_out(gen8_out));
assign random_out = gen1_out  ^ gen2_out;// ^ gen3_out ^ gen4_out ^ gen5_out ^ gen6_out ^ gen7_out ^ gen8_out;
//tutaj w zależności od dodatkowego parametru dajemy różne wyjścia:

//SHA3 
sha3 sha3_(
           .clk(clk),
           .nreset(reset),
           .w(sha3_we),
           .addr(sha3_address),
           .din(sha3_din),
           .dout(sha3_dout),
           .init(sha3_init),
           .next(sha3_next),
           .ready(sha3_ready)
           );

//module sha3(    input wire          clk,
//                input wire 	     nreset,
//                input wire 	     w,
//                input wire [ 8:2]    addr,
//                input wire [32-1:0]  din,
//                output wire [32-1:0] dout,
//                input wire 	     init,
//                input wire 	     next,
//                output wire 	     ready);

assign writed_words_counter_wire = writed_words_counter;

//STATE MACHINE
always @(posedge clk)
begin
    if(reset)
        begin
        state = starting;
        generated_bits_counter = 16'h0000;
        generating_hash_counter = 0;
        digest_data = 0;
        random_bits = 0;
        writed_words_counter = 0;
        readed_words_counter = 0;
        end
    else
    begin
    case(state)
        starting: begin
            state <= generating;
        end
        
        generating: begin
            if(generated_bits_counter < CHUNK_SIZE)
            begin
                random_bits[generated_bits_counter] <= random_out;
                generated_bits_counter <= generated_bits_counter + 1;
            end
            if(generated_bits_counter == CHUNK_SIZE)
            begin
                state <= generated;
                generated_bits_counter <= 16'h0000; 
            end
         end
         
         generated: begin
            state <= writing_to_sha;
         end
         
         writing_to_sha: begin//zapisywanie danych do sha po 32 bity ///3
            case(writed_words_counter[5:0])
                6'b000000 : sha3_address <= ADDR_BLOCK0;
                6'b000001 : sha3_address <= ADDR_BLOCK1;
                6'b000010 : sha3_address <= ADDR_BLOCK2;
                6'b000011 : sha3_address <= ADDR_BLOCK3;
                6'b000100 : sha3_address <= ADDR_BLOCK4;
                6'b000101 : sha3_address <= ADDR_BLOCK5;
                6'b000110 : sha3_address <= ADDR_BLOCK6;
                6'b000111 : sha3_address <= ADDR_BLOCK7;
                6'b001000 : sha3_address <= ADDR_BLOCK8;
                6'b001001 : sha3_address <= ADDR_BLOCK9;
                6'b001010 : sha3_address <= ADDR_BLOCK10;
                6'b001011 : sha3_address <= ADDR_BLOCK11;
                6'b001100 : sha3_address <= ADDR_BLOCK12;
                6'b001101 : sha3_address <= ADDR_BLOCK13;
                6'b001110 : sha3_address <= ADDR_BLOCK14;
                6'b001111 : sha3_address <= ADDR_BLOCK15;
                6'b010000 : sha3_address <= ADDR_BLOCK16;
                6'b010001 : sha3_address <= ADDR_BLOCK17;
                6'b010010 : sha3_address <= ADDR_BLOCK18;
                6'b010011 : sha3_address <= ADDR_BLOCK19;
                6'b010100 : sha3_address <= ADDR_BLOCK20;
                6'b010101 : sha3_address <= ADDR_BLOCK21;
                6'b010110 : sha3_address <= ADDR_BLOCK22;
                6'b010111 : sha3_address <= ADDR_BLOCK23;
                6'b011000 : sha3_address <= ADDR_BLOCK24;
                6'b011001 : sha3_address <= ADDR_BLOCK25;
                6'b011010 : sha3_address <= ADDR_BLOCK26;
                6'b011011 : sha3_address <= ADDR_BLOCK27;
                6'b011100 : sha3_address <= ADDR_BLOCK28;
                6'b011101 : sha3_address <= ADDR_BLOCK29;
                6'b011110 : sha3_address <= ADDR_BLOCK30;
                6'b011111 : sha3_address <= ADDR_BLOCK31;
                6'b100000 : sha3_address <= ADDR_BLOCK32;
                6'b100001 : sha3_address <= ADDR_BLOCK33;
                6'b100010 : sha3_address <= ADDR_BLOCK34;
                6'b100011 : sha3_address <= ADDR_BLOCK35;
                6'b100100 : sha3_address <= ADDR_BLOCK36;
                6'b100101 : sha3_address <= ADDR_BLOCK37;
                6'b100110 : sha3_address <= ADDR_BLOCK38;
                6'b100111 : sha3_address <= ADDR_BLOCK39;
                6'b101000 : sha3_address <= ADDR_BLOCK40;
                6'b101001 : sha3_address <= ADDR_BLOCK41;
                6'b101010 : sha3_address <= ADDR_BLOCK42;
                6'b101011 : sha3_address <= ADDR_BLOCK43;
                6'b101100 : sha3_address <= ADDR_BLOCK44;
                6'b101101 : sha3_address <= ADDR_BLOCK45;
                6'b101110 : sha3_address <= ADDR_BLOCK46;
                6'b101111 : sha3_address <= ADDR_BLOCK47;
                6'b110000 : sha3_address <= ADDR_BLOCK48;
                6'b110001 : sha3_address <= ADDR_BLOCK49;
                default : sha3_address <= ADDR_BLOCK0;
            endcase 
            
            case(writed_words_counter)
                10'h000 :  sha3_din <= random_bits[31:0];
                10'h001 :  sha3_din <= random_bits[63:32];
                10'h002 :  sha3_din <= random_bits[95:64];
                10'h003 :  sha3_din <= random_bits[127:96];
                10'h004 :  sha3_din <= random_bits[159:128];
                10'h005 :  sha3_din <= random_bits[191:160];
                10'h006 :  sha3_din <= random_bits[223:192];
                10'h007 :  sha3_din <= random_bits[255:224];
                10'h008 :  sha3_din <= random_bits[287:256];
                10'h009 :  sha3_din <= random_bits[319:288];
                10'h00a :  sha3_din <= random_bits[351:320];
                10'h00b :  sha3_din <= random_bits[383:352];
                10'h00c :  sha3_din <= random_bits[415:384];
                10'h00d :  sha3_din <= random_bits[447:416];
                10'h00e :  sha3_din <= random_bits[479:448];
                10'h00f :  sha3_din <= random_bits[511:480];
                10'h010 :  sha3_din <= random_bits[543:512];
                10'h011 :  sha3_din <= random_bits[575:544];
                10'h012 :  sha3_din <= random_bits[607:576];
                10'h013 :  sha3_din <= random_bits[639:608];
                10'h014 :  sha3_din <= random_bits[671:640];
                10'h015 :  sha3_din <= random_bits[703:672];
                10'h016 :  sha3_din <= random_bits[735:704];
                10'h017 :  sha3_din <= random_bits[767:736];
                10'h018 :  sha3_din <= random_bits[799:768];
                10'h019 :  sha3_din <= random_bits[831:800];
                10'h01a :  sha3_din <= random_bits[863:832];
                10'h01b :  sha3_din <= random_bits[895:864];
                10'h01c :  sha3_din <= random_bits[927:896];
                10'h01d :  sha3_din <= random_bits[959:928];
                10'h01e :  sha3_din <= random_bits[991:960];
                10'h01f :  sha3_din <= random_bits[1023:992];
                // 10'h020 :  sha3_din <= random_bits[1055:1024];
                // 10'h021 :  sha3_din <= random_bits[1087:1056];
                // 10'h022 :  sha3_din <= random_bits[1119:1088];
                // 10'h023 :  sha3_din <= random_bits[1151:1120];
                // 10'h024 :  sha3_din <= random_bits[1183:1152];
                // 10'h025 :  sha3_din <= random_bits[1215:1184];
                // 10'h026 :  sha3_din <= random_bits[1247:1216];
                // 10'h027 :  sha3_din <= random_bits[1279:1248];
                // 10'h028 :  sha3_din <= random_bits[1311:1280];
                // 10'h029 :  sha3_din <= random_bits[1343:1312];
                // 10'h02a :  sha3_din <= random_bits[1375:1344];
                // 10'h02b :  sha3_din <= random_bits[1407:1376];
                // 10'h02c :  sha3_din <= random_bits[1439:1408];
                // 10'h02d :  sha3_din <= random_bits[1471:1440];
                // 10'h02e :  sha3_din <= random_bits[1503:1472];
                // 10'h02f :  sha3_din <= random_bits[1535:1504];
                // 10'h030 :  sha3_din <= random_bits[1567:1536];
                // 10'h031 :  sha3_din <= random_bits[1599:1568];
                // 10'h032 :  sha3_din <= random_bits[1631:1600];
                // 10'h033 :  sha3_din <= random_bits[1663:1632];
                // 10'h034 :  sha3_din <= random_bits[1695:1664];
                // 10'h035 :  sha3_din <= random_bits[1727:1696];
                // 10'h036 :  sha3_din <= random_bits[1759:1728];
                // 10'h037 :  sha3_din <= random_bits[1791:1760];
                // 10'h038 :  sha3_din <= random_bits[1823:1792];
                // 10'h039 :  sha3_din <= random_bits[1855:1824];
                // 10'h03a :  sha3_din <= random_bits[1887:1856];
                // 10'h03b :  sha3_din <= random_bits[1919:1888];
                // 10'h03c :  sha3_din <= random_bits[1951:1920];
                // 10'h03d :  sha3_din <= random_bits[1983:1952];
                // 10'h03e :  sha3_din <= random_bits[2015:1984];
                // 10'h03f :  sha3_din <= random_bits[2047:2016];
                // 10'h040 :  sha3_din <= random_bits[2079:2048];
                // 10'h041 :  sha3_din <= random_bits[2111:2080];
                // 10'h042 :  sha3_din <= random_bits[2143:2112];
                // 10'h043 :  sha3_din <= random_bits[2175:2144];
                // 10'h044 :  sha3_din <= random_bits[2207:2176];
                // 10'h045 :  sha3_din <= random_bits[2239:2208];
                // 10'h046 :  sha3_din <= random_bits[2271:2240];
                // 10'h047 :  sha3_din <= random_bits[2303:2272];
                // 10'h048 :  sha3_din <= random_bits[2335:2304];
                // 10'h049 :  sha3_din <= random_bits[2367:2336];
                // 10'h04a :  sha3_din <= random_bits[2399:2368];
                // 10'h04b :  sha3_din <= random_bits[2431:2400];
                // 10'h04c :  sha3_din <= random_bits[2463:2432];
                // 10'h04d :  sha3_din <= random_bits[2495:2464];
                // 10'h04e :  sha3_din <= random_bits[2527:2496];
                // 10'h04f :  sha3_din <= random_bits[2559:2528];
                // 10'h050 :  sha3_din <= random_bits[2591:2560];
                // 10'h051 :  sha3_din <= random_bits[2623:2592];
                // 10'h052 :  sha3_din <= random_bits[2655:2624];
                // 10'h053 :  sha3_din <= random_bits[2687:2656];
                // 10'h054 :  sha3_din <= random_bits[2719:2688];
                // 10'h055 :  sha3_din <= random_bits[2751:2720];
                // 10'h056 :  sha3_din <= random_bits[2783:2752];
                // 10'h057 :  sha3_din <= random_bits[2815:2784];
                // 10'h058 :  sha3_din <= random_bits[2847:2816];
                // 10'h059 :  sha3_din <= random_bits[2879:2848];
                // 10'h05a :  sha3_din <= random_bits[2911:2880];
                // 10'h05b :  sha3_din <= random_bits[2943:2912];
                // 10'h05c :  sha3_din <= random_bits[2975:2944];
                // 10'h05d :  sha3_din <= random_bits[3007:2976];
                // 10'h05e :  sha3_din <= random_bits[3039:3008];
                // 10'h05f :  sha3_din <= random_bits[3071:3040];
                // 10'h060 :  sha3_din <= random_bits[3103:3072];
                // 10'h061 :  sha3_din <= random_bits[3135:3104];
                // 10'h062 :  sha3_din <= random_bits[3167:3136];
                // 10'h063 :  sha3_din <= random_bits[3199:3168];
                // 10'h064 :  sha3_din <= random_bits[3231:3200];
                // 10'h065 :  sha3_din <= random_bits[3263:3232];
                // 10'h066 :  sha3_din <= random_bits[3295:3264];
                // 10'h067 :  sha3_din <= random_bits[3327:3296];
                // 10'h068 :  sha3_din <= random_bits[3359:3328];
                // 10'h069 :  sha3_din <= random_bits[3391:3360];
                // 10'h06a :  sha3_din <= random_bits[3423:3392];
                // 10'h06b :  sha3_din <= random_bits[3455:3424];
                // 10'h06c :  sha3_din <= random_bits[3487:3456];
                // 10'h06d :  sha3_din <= random_bits[3519:3488];
                // 10'h06e :  sha3_din <= random_bits[3551:3520];
                // 10'h06f :  sha3_din <= random_bits[3583:3552];
                // 10'h070 :  sha3_din <= random_bits[3615:3584];
                // 10'h071 :  sha3_din <= random_bits[3647:3616];
                // 10'h072 :  sha3_din <= random_bits[3679:3648];
                // 10'h073 :  sha3_din <= random_bits[3711:3680];
                // 10'h074 :  sha3_din <= random_bits[3743:3712];
                // 10'h075 :  sha3_din <= random_bits[3775:3744];
                // 10'h076 :  sha3_din <= random_bits[3807:3776];
                // 10'h077 :  sha3_din <= random_bits[3839:3808];
                // 10'h078 :  sha3_din <= random_bits[3871:3840];
                // 10'h079 :  sha3_din <= random_bits[3903:3872];
                // 10'h07a :  sha3_din <= random_bits[3935:3904];
                // 10'h07b :  sha3_din <= random_bits[3967:3936];
                // 10'h07c :  sha3_din <= random_bits[3999:3968];
                // 10'h07d :  sha3_din <= random_bits[4031:4000];
                // 10'h07e :  sha3_din <= random_bits[4063:4032];
                // 10'h07f :  sha3_din <= random_bits[4095:4064];
                // 10'h080 :  sha3_din <= random_bits[4127:4096];
                // 10'h081 :  sha3_din <= random_bits[4159:4128];
                // 10'h082 :  sha3_din <= random_bits[4191:4160];
                // 10'h083 :  sha3_din <= random_bits[4223:4192];
                // 10'h084 :  sha3_din <= random_bits[4255:4224];
                // 10'h085 :  sha3_din <= random_bits[4287:4256];
                // 10'h086 :  sha3_din <= random_bits[4319:4288];
                // 10'h087 :  sha3_din <= random_bits[4351:4320];
                // 10'h088 :  sha3_din <= random_bits[4383:4352];
                // 10'h089 :  sha3_din <= random_bits[4415:4384];
                // 10'h08a :  sha3_din <= random_bits[4447:4416];
                // 10'h08b :  sha3_din <= random_bits[4479:4448];
                // 10'h08c :  sha3_din <= random_bits[4511:4480];
                // 10'h08d :  sha3_din <= random_bits[4543:4512];
                // 10'h08e :  sha3_din <= random_bits[4575:4544];
                // 10'h08f :  sha3_din <= random_bits[4607:4576];
                // 10'h090 :  sha3_din <= random_bits[4639:4608];
                // 10'h091 :  sha3_din <= random_bits[4671:4640];
                // 10'h092 :  sha3_din <= random_bits[4703:4672];
                // 10'h093 :  sha3_din <= random_bits[4735:4704];
                // 10'h094 :  sha3_din <= random_bits[4767:4736];
                // 10'h095 :  sha3_din <= random_bits[4799:4768];
                // 10'h096 :  sha3_din <= random_bits[4831:4800];
                // 10'h097 :  sha3_din <= random_bits[4863:4832];
                // 10'h098 :  sha3_din <= random_bits[4895:4864];
                // 10'h099 :  sha3_din <= random_bits[4927:4896];
                // 10'h09a :  sha3_din <= random_bits[4959:4928];
                // 10'h09b :  sha3_din <= random_bits[4991:4960];
                // 10'h09c :  sha3_din <= random_bits[5023:4992];
                // 10'h09d :  sha3_din <= random_bits[5055:5024];
                // 10'h09e :  sha3_din <= random_bits[5087:5056];
                // 10'h09f :  sha3_din <= random_bits[5119:5088];
                // 10'h0a0 :  sha3_din <= random_bits[5151:5120];
                // 10'h0a1 :  sha3_din <= random_bits[5183:5152];
                // 10'h0a2 :  sha3_din <= random_bits[5215:5184];
                // 10'h0a3 :  sha3_din <= random_bits[5247:5216];
                // 10'h0a4 :  sha3_din <= random_bits[5279:5248];
                // 10'h0a5 :  sha3_din <= random_bits[5311:5280];
                // 10'h0a6 :  sha3_din <= random_bits[5343:5312];
                // 10'h0a7 :  sha3_din <= random_bits[5375:5344];
                // 10'h0a8 :  sha3_din <= random_bits[5407:5376];
                // 10'h0a9 :  sha3_din <= random_bits[5439:5408];
                // 10'h0aa :  sha3_din <= random_bits[5471:5440];
                // 10'h0ab :  sha3_din <= random_bits[5503:5472];
                // 10'h0ac :  sha3_din <= random_bits[5535:5504];
                // 10'h0ad :  sha3_din <= random_bits[5567:5536];
                // 10'h0ae :  sha3_din <= random_bits[5599:5568];
                // 10'h0af :  sha3_din <= random_bits[5631:5600];
                // 10'h0b0 :  sha3_din <= random_bits[5663:5632];
                // 10'h0b1 :  sha3_din <= random_bits[5695:5664];
                // 10'h0b2 :  sha3_din <= random_bits[5727:5696];
                // 10'h0b3 :  sha3_din <= random_bits[5759:5728];
                // 10'h0b4 :  sha3_din <= random_bits[5791:5760];
                // 10'h0b5 :  sha3_din <= random_bits[5823:5792];
                // 10'h0b6 :  sha3_din <= random_bits[5855:5824];
                // 10'h0b7 :  sha3_din <= random_bits[5887:5856];
                // 10'h0b8 :  sha3_din <= random_bits[5919:5888];
                // 10'h0b9 :  sha3_din <= random_bits[5951:5920];
                // 10'h0ba :  sha3_din <= random_bits[5983:5952];
                // 10'h0bb :  sha3_din <= random_bits[6015:5984];
                // 10'h0bc :  sha3_din <= random_bits[6047:6016];
                // 10'h0bd :  sha3_din <= random_bits[6079:6048];
                // 10'h0be :  sha3_din <= random_bits[6111:6080];
                // 10'h0bf :  sha3_din <= random_bits[6143:6112];
                // 10'h0c0 :  sha3_din <= random_bits[6175:6144];
                // 10'h0c1 :  sha3_din <= random_bits[6207:6176];
                // 10'h0c2 :  sha3_din <= random_bits[6239:6208];
                // 10'h0c3 :  sha3_din <= random_bits[6271:6240];
                // 10'h0c4 :  sha3_din <= random_bits[6303:6272];
                // 10'h0c5 :  sha3_din <= random_bits[6335:6304];
                // 10'h0c6 :  sha3_din <= random_bits[6367:6336];
                // 10'h0c7 :  sha3_din <= random_bits[6399:6368];
                // 10'h0c8 :  sha3_din <= random_bits[6431:6400];
                // 10'h0c9 :  sha3_din <= random_bits[6463:6432];
                // 10'h0ca :  sha3_din <= random_bits[6495:6464];
                // 10'h0cb :  sha3_din <= random_bits[6527:6496];
                // 10'h0cc :  sha3_din <= random_bits[6559:6528];
                // 10'h0cd :  sha3_din <= random_bits[6591:6560];
                // 10'h0ce :  sha3_din <= random_bits[6623:6592];
                // 10'h0cf :  sha3_din <= random_bits[6655:6624];
                // 10'h0d0 :  sha3_din <= random_bits[6687:6656];
                // 10'h0d1 :  sha3_din <= random_bits[6719:6688];
                // 10'h0d2 :  sha3_din <= random_bits[6751:6720];
                // 10'h0d3 :  sha3_din <= random_bits[6783:6752];
                // 10'h0d4 :  sha3_din <= random_bits[6815:6784];
                // 10'h0d5 :  sha3_din <= random_bits[6847:6816];
                // 10'h0d6 :  sha3_din <= random_bits[6879:6848];
                // 10'h0d7 :  sha3_din <= random_bits[6911:6880];
                // 10'h0d8 :  sha3_din <= random_bits[6943:6912];
                // 10'h0d9 :  sha3_din <= random_bits[6975:6944];
                // 10'h0da :  sha3_din <= random_bits[7007:6976];
                // 10'h0db :  sha3_din <= random_bits[7039:7008];
                // 10'h0dc :  sha3_din <= random_bits[7071:7040];
                // 10'h0dd :  sha3_din <= random_bits[7103:7072];
                // 10'h0de :  sha3_din <= random_bits[7135:7104];
                // 10'h0df :  sha3_din <= random_bits[7167:7136];
                // 10'h0e0 :  sha3_din <= random_bits[7199:7168];
                // 10'h0e1 :  sha3_din <= random_bits[7231:7200];
                // 10'h0e2 :  sha3_din <= random_bits[7263:7232];
                // 10'h0e3 :  sha3_din <= random_bits[7295:7264];
                // 10'h0e4 :  sha3_din <= random_bits[7327:7296];
                // 10'h0e5 :  sha3_din <= random_bits[7359:7328];
                // 10'h0e6 :  sha3_din <= random_bits[7391:7360];
                // 10'h0e7 :  sha3_din <= random_bits[7423:7392];
                // 10'h0e8 :  sha3_din <= random_bits[7455:7424];
                // 10'h0e9 :  sha3_din <= random_bits[7487:7456];
                // 10'h0ea :  sha3_din <= random_bits[7519:7488];
                // 10'h0eb :  sha3_din <= random_bits[7551:7520];
                // 10'h0ec :  sha3_din <= random_bits[7583:7552];
                // 10'h0ed :  sha3_din <= random_bits[7615:7584];
                // 10'h0ee :  sha3_din <= random_bits[7647:7616];
                // 10'h0ef :  sha3_din <= random_bits[7679:7648];
                // 10'h0f0 :  sha3_din <= random_bits[7711:7680];
                // 10'h0f1 :  sha3_din <= random_bits[7743:7712];
                // 10'h0f2 :  sha3_din <= random_bits[7775:7744];
                // 10'h0f3 :  sha3_din <= random_bits[7807:7776];
                // 10'h0f4 :  sha3_din <= random_bits[7839:7808];
                // 10'h0f5 :  sha3_din <= random_bits[7871:7840];
                // 10'h0f6 :  sha3_din <= random_bits[7903:7872];
                // 10'h0f7 :  sha3_din <= random_bits[7935:7904];
                // 10'h0f8 :  sha3_din <= random_bits[7967:7936];
                // 10'h0f9 :  sha3_din <= random_bits[7999:7968];
                // 10'h0fa :  sha3_din <= random_bits[8031:8000];
                // 10'h0fb :  sha3_din <= random_bits[8063:8032];
                // 10'h0fc :  sha3_din <= random_bits[8095:8064];
                // 10'h0fd :  sha3_din <= random_bits[8127:8096];
                // 10'h0fe :  sha3_din <= random_bits[8159:8128];
                // 10'h0ff :  sha3_din <= random_bits[8191:8160];
                // 10'h100 :  sha3_din <= random_bits[8223:8192];
                // 10'h101 :  sha3_din <= random_bits[8255:8224];
                // 10'h102 :  sha3_din <= random_bits[8287:8256];
                // 10'h103 :  sha3_din <= random_bits[8319:8288];
                // 10'h104 :  sha3_din <= random_bits[8351:8320];
                // 10'h105 :  sha3_din <= random_bits[8383:8352];
                // 10'h106 :  sha3_din <= random_bits[8415:8384];
                // 10'h107 :  sha3_din <= random_bits[8447:8416];
                // 10'h108 :  sha3_din <= random_bits[8479:8448];
                // 10'h109 :  sha3_din <= random_bits[8511:8480];
                // 10'h10a :  sha3_din <= random_bits[8543:8512];
                // 10'h10b :  sha3_din <= random_bits[8575:8544];
                // 10'h10c :  sha3_din <= random_bits[8607:8576];
                // 10'h10d :  sha3_din <= random_bits[8639:8608];
                // 10'h10e :  sha3_din <= random_bits[8671:8640];
                // 10'h10f :  sha3_din <= random_bits[8703:8672];
                // 10'h110 :  sha3_din <= random_bits[8735:8704];
                // 10'h111 :  sha3_din <= random_bits[8767:8736];
                // 10'h112 :  sha3_din <= random_bits[8799:8768];
                // 10'h113 :  sha3_din <= random_bits[8831:8800];
                // 10'h114 :  sha3_din <= random_bits[8863:8832];
                // 10'h115 :  sha3_din <= random_bits[8895:8864];
                // 10'h116 :  sha3_din <= random_bits[8927:8896];
                // 10'h117 :  sha3_din <= random_bits[8959:8928];
                // 10'h118 :  sha3_din <= random_bits[8991:8960];
                // 10'h119 :  sha3_din <= random_bits[9023:8992];
                // 10'h11a :  sha3_din <= random_bits[9055:9024];
                // 10'h11b :  sha3_din <= random_bits[9087:9056];
                // 10'h11c :  sha3_din <= random_bits[9119:9088];
                // 10'h11d :  sha3_din <= random_bits[9151:9120];
                // 10'h11e :  sha3_din <= random_bits[9183:9152];
                // 10'h11f :  sha3_din <= random_bits[9215:9184];
                // 10'h120 :  sha3_din <= random_bits[9247:9216];
                // 10'h121 :  sha3_din <= random_bits[9279:9248];
                // 10'h122 :  sha3_din <= random_bits[9311:9280];
                // 10'h123 :  sha3_din <= random_bits[9343:9312];
                // 10'h124 :  sha3_din <= random_bits[9375:9344];
                // 10'h125 :  sha3_din <= random_bits[9407:9376];
                // 10'h126 :  sha3_din <= random_bits[9439:9408];
                // 10'h127 :  sha3_din <= random_bits[9471:9440];
                // 10'h128 :  sha3_din <= random_bits[9503:9472];
                // 10'h129 :  sha3_din <= random_bits[9535:9504];
                // 10'h12a :  sha3_din <= random_bits[9567:9536];
                // 10'h12b :  sha3_din <= random_bits[9599:9568];
                // 10'h12c :  sha3_din <= random_bits[9631:9600];
                // 10'h12d :  sha3_din <= random_bits[9663:9632];
                // 10'h12e :  sha3_din <= random_bits[9695:9664];
                // 10'h12f :  sha3_din <= random_bits[9727:9696];
                // 10'h130 :  sha3_din <= random_bits[9759:9728];
                // 10'h131 :  sha3_din <= random_bits[9791:9760];
                // 10'h132 :  sha3_din <= random_bits[9823:9792];
                // 10'h133 :  sha3_din <= random_bits[9855:9824];
                // 10'h134 :  sha3_din <= random_bits[9887:9856];
                // 10'h135 :  sha3_din <= random_bits[9919:9888];
                // 10'h136 :  sha3_din <= random_bits[9951:9920];
                // 10'h137 :  sha3_din <= random_bits[9983:9952];
                // 10'h138 :  sha3_din <= random_bits[10015:9984];
                // 10'h139 :  sha3_din <= random_bits[10047:10016];
                // 10'h13a :  sha3_din <= random_bits[10079:10048];
                // 10'h13b :  sha3_din <= random_bits[10111:10080];
                // 10'h13c :  sha3_din <= random_bits[10143:10112];
                // 10'h13d :  sha3_din <= random_bits[10175:10144];
                // 10'h13e :  sha3_din <= random_bits[10207:10176];
                // 10'h13f :  sha3_din <= random_bits[10239:10208];
                // 10'h140 :  sha3_din <= random_bits[10271:10240];
                // 10'h141 :  sha3_din <= random_bits[10303:10272];
                // 10'h142 :  sha3_din <= random_bits[10335:10304];
                // 10'h143 :  sha3_din <= random_bits[10367:10336];
                // 10'h144 :  sha3_din <= random_bits[10399:10368];
                // 10'h145 :  sha3_din <= random_bits[10431:10400];
                // 10'h146 :  sha3_din <= random_bits[10463:10432];
                // 10'h147 :  sha3_din <= random_bits[10495:10464];
                // 10'h148 :  sha3_din <= random_bits[10527:10496];
                // 10'h149 :  sha3_din <= random_bits[10559:10528];
                // 10'h14a :  sha3_din <= random_bits[10591:10560];
                // 10'h14b :  sha3_din <= random_bits[10623:10592];
                // 10'h14c :  sha3_din <= random_bits[10655:10624];
                // 10'h14d :  sha3_din <= random_bits[10687:10656];
                // 10'h14e :  sha3_din <= random_bits[10719:10688];
                // 10'h14f :  sha3_din <= random_bits[10751:10720];
                // 10'h150 :  sha3_din <= random_bits[10783:10752];
                // 10'h151 :  sha3_din <= random_bits[10815:10784];
                // 10'h152 :  sha3_din <= random_bits[10847:10816];
                // 10'h153 :  sha3_din <= random_bits[10879:10848];
                // 10'h154 :  sha3_din <= random_bits[10911:10880];
                // 10'h155 :  sha3_din <= random_bits[10943:10912];
                // 10'h156 :  sha3_din <= random_bits[10975:10944];
                // 10'h157 :  sha3_din <= random_bits[11007:10976];
                // 10'h158 :  sha3_din <= random_bits[11039:11008];
                // 10'h159 :  sha3_din <= random_bits[11071:11040];
                // 10'h15a :  sha3_din <= random_bits[11103:11072];
                // 10'h15b :  sha3_din <= random_bits[11135:11104];
                // 10'h15c :  sha3_din <= random_bits[11167:11136];
                // 10'h15d :  sha3_din <= random_bits[11199:11168];
                // 10'h15e :  sha3_din <= random_bits[11231:11200];
                // 10'h15f :  sha3_din <= random_bits[11263:11232];
                // 10'h160 :  sha3_din <= random_bits[11295:11264];
                // 10'h161 :  sha3_din <= random_bits[11327:11296];
                // 10'h162 :  sha3_din <= random_bits[11359:11328];
                // 10'h163 :  sha3_din <= random_bits[11391:11360];
                // 10'h164 :  sha3_din <= random_bits[11423:11392];
                // 10'h165 :  sha3_din <= random_bits[11455:11424];
                // 10'h166 :  sha3_din <= random_bits[11487:11456];
                // 10'h167 :  sha3_din <= random_bits[11519:11488];
                // 10'h168 :  sha3_din <= random_bits[11551:11520];
                // 10'h169 :  sha3_din <= random_bits[11583:11552];
                // 10'h16a :  sha3_din <= random_bits[11615:11584];
                // 10'h16b :  sha3_din <= random_bits[11647:11616];
                // 10'h16c :  sha3_din <= random_bits[11679:11648];
                // 10'h16d :  sha3_din <= random_bits[11711:11680];
                // 10'h16e :  sha3_din <= random_bits[11743:11712];
                // 10'h16f :  sha3_din <= random_bits[11775:11744];
                // 10'h170 :  sha3_din <= random_bits[11807:11776];
                // 10'h171 :  sha3_din <= random_bits[11839:11808];
                // 10'h172 :  sha3_din <= random_bits[11871:11840];
                // 10'h173 :  sha3_din <= random_bits[11903:11872];
                // 10'h174 :  sha3_din <= random_bits[11935:11904];
                // 10'h175 :  sha3_din <= random_bits[11967:11936];
                // 10'h176 :  sha3_din <= random_bits[11999:11968];
                // 10'h177 :  sha3_din <= random_bits[12031:12000];
                // 10'h178 :  sha3_din <= random_bits[12063:12032];
                // 10'h179 :  sha3_din <= random_bits[12095:12064];
                // 10'h17a :  sha3_din <= random_bits[12127:12096];
                // 10'h17b :  sha3_din <= random_bits[12159:12128];
                // 10'h17c :  sha3_din <= random_bits[12191:12160];
                // 10'h17d :  sha3_din <= random_bits[12223:12192];
                // 10'h17e :  sha3_din <= random_bits[12255:12224];
                // 10'h17f :  sha3_din <= random_bits[12287:12256];
                // 10'h180 :  sha3_din <= random_bits[12319:12288];
                // 10'h181 :  sha3_din <= random_bits[12351:12320];
                // 10'h182 :  sha3_din <= random_bits[12383:12352];
                // 10'h183 :  sha3_din <= random_bits[12415:12384];
                // 10'h184 :  sha3_din <= random_bits[12447:12416];
                // 10'h185 :  sha3_din <= random_bits[12479:12448];
                // 10'h186 :  sha3_din <= random_bits[12511:12480];
                // 10'h187 :  sha3_din <= random_bits[12543:12512];
                // 10'h188 :  sha3_din <= random_bits[12575:12544];
                // 10'h189 :  sha3_din <= random_bits[12607:12576];
                // 10'h18a :  sha3_din <= random_bits[12639:12608];
                // 10'h18b :  sha3_din <= random_bits[12671:12640];
                // 10'h18c :  sha3_din <= random_bits[12703:12672];
                // 10'h18d :  sha3_din <= random_bits[12735:12704];
                // 10'h18e :  sha3_din <= random_bits[12767:12736];
                // 10'h18f :  sha3_din <= random_bits[12799:12768];
                // 10'h190 :  sha3_din <= random_bits[12831:12800];
                // 10'h191 :  sha3_din <= random_bits[12863:12832];
                // 10'h192 :  sha3_din <= random_bits[12895:12864];
                // 10'h193 :  sha3_din <= random_bits[12927:12896];
                // 10'h194 :  sha3_din <= random_bits[12959:12928];
                // 10'h195 :  sha3_din <= random_bits[12991:12960];
                // 10'h196 :  sha3_din <= random_bits[13023:12992];
                // 10'h197 :  sha3_din <= random_bits[13055:13024];
                // 10'h198 :  sha3_din <= random_bits[13087:13056];
                // 10'h199 :  sha3_din <= random_bits[13119:13088];
                // 10'h19a :  sha3_din <= random_bits[13151:13120];
                // 10'h19b :  sha3_din <= random_bits[13183:13152];
                // 10'h19c :  sha3_din <= random_bits[13215:13184];
                // 10'h19d :  sha3_din <= random_bits[13247:13216];
                // 10'h19e :  sha3_din <= random_bits[13279:13248];
                // 10'h19f :  sha3_din <= random_bits[13311:13280];
                // 10'h1a0 :  sha3_din <= random_bits[13343:13312];
                // 10'h1a1 :  sha3_din <= random_bits[13375:13344];
                // 10'h1a2 :  sha3_din <= random_bits[13407:13376];
                // 10'h1a3 :  sha3_din <= random_bits[13439:13408];
                // 10'h1a4 :  sha3_din <= random_bits[13471:13440];
                // 10'h1a5 :  sha3_din <= random_bits[13503:13472];
                // 10'h1a6 :  sha3_din <= random_bits[13535:13504];
                // 10'h1a7 :  sha3_din <= random_bits[13567:13536];
                // 10'h1a8 :  sha3_din <= random_bits[13599:13568];
                // 10'h1a9 :  sha3_din <= random_bits[13631:13600];
                // 10'h1aa :  sha3_din <= random_bits[13663:13632];
                // 10'h1ab :  sha3_din <= random_bits[13695:13664];
                // 10'h1ac :  sha3_din <= random_bits[13727:13696];
                // 10'h1ad :  sha3_din <= random_bits[13759:13728];
                // 10'h1ae :  sha3_din <= random_bits[13791:13760];
                // 10'h1af :  sha3_din <= random_bits[13823:13792];
                // 10'h1b0 :  sha3_din <= random_bits[13855:13824];
                // 10'h1b1 :  sha3_din <= random_bits[13887:13856];
                // 10'h1b2 :  sha3_din <= random_bits[13919:13888];
                // 10'h1b3 :  sha3_din <= random_bits[13951:13920];
                // 10'h1b4 :  sha3_din <= random_bits[13983:13952];
                // 10'h1b5 :  sha3_din <= random_bits[14015:13984];
                // 10'h1b6 :  sha3_din <= random_bits[14047:14016];
                // 10'h1b7 :  sha3_din <= random_bits[14079:14048];
                // 10'h1b8 :  sha3_din <= random_bits[14111:14080];
                // 10'h1b9 :  sha3_din <= random_bits[14143:14112];
                // 10'h1ba :  sha3_din <= random_bits[14175:14144];
                // 10'h1bb :  sha3_din <= random_bits[14207:14176];
                // 10'h1bc :  sha3_din <= random_bits[14239:14208];
                // 10'h1bd :  sha3_din <= random_bits[14271:14240];
                // 10'h1be :  sha3_din <= random_bits[14303:14272];
                // 10'h1bf :  sha3_din <= random_bits[14335:14304];
                // 10'h1c0 :  sha3_din <= random_bits[14367:14336];
                // 10'h1c1 :  sha3_din <= random_bits[14399:14368];
                // 10'h1c2 :  sha3_din <= random_bits[14431:14400];
                // 10'h1c3 :  sha3_din <= random_bits[14463:14432];
                // 10'h1c4 :  sha3_din <= random_bits[14495:14464];
                // 10'h1c5 :  sha3_din <= random_bits[14527:14496];
                // 10'h1c6 :  sha3_din <= random_bits[14559:14528];
                // 10'h1c7 :  sha3_din <= random_bits[14591:14560];
                // 10'h1c8 :  sha3_din <= random_bits[14623:14592];
                // 10'h1c9 :  sha3_din <= random_bits[14655:14624];
                // 10'h1ca :  sha3_din <= random_bits[14687:14656];
                // 10'h1cb :  sha3_din <= random_bits[14719:14688];
                // 10'h1cc :  sha3_din <= random_bits[14751:14720];
                // 10'h1cd :  sha3_din <= random_bits[14783:14752];
                // 10'h1ce :  sha3_din <= random_bits[14815:14784];
                // 10'h1cf :  sha3_din <= random_bits[14847:14816];
                // 10'h1d0 :  sha3_din <= random_bits[14879:14848];
                // 10'h1d1 :  sha3_din <= random_bits[14911:14880];
                // 10'h1d2 :  sha3_din <= random_bits[14943:14912];
                // 10'h1d3 :  sha3_din <= random_bits[14975:14944];
                // 10'h1d4 :  sha3_din <= random_bits[15007:14976];
                // 10'h1d5 :  sha3_din <= random_bits[15039:15008];
                // 10'h1d6 :  sha3_din <= random_bits[15071:15040];
                // 10'h1d7 :  sha3_din <= random_bits[15103:15072];
                // 10'h1d8 :  sha3_din <= random_bits[15135:15104];
                // 10'h1d9 :  sha3_din <= random_bits[15167:15136];
                // 10'h1da :  sha3_din <= random_bits[15199:15168];
                // 10'h1db :  sha3_din <= random_bits[15231:15200];
                // 10'h1dc :  sha3_din <= random_bits[15263:15232];
                // 10'h1dd :  sha3_din <= random_bits[15295:15264];
                // 10'h1de :  sha3_din <= random_bits[15327:15296];
                // 10'h1df :  sha3_din <= random_bits[15359:15328];
                // 10'h1e0 :  sha3_din <= random_bits[15391:15360];
                // 10'h1e1 :  sha3_din <= random_bits[15423:15392];
                // 10'h1e2 :  sha3_din <= random_bits[15455:15424];
                // 10'h1e3 :  sha3_din <= random_bits[15487:15456];
                // 10'h1e4 :  sha3_din <= random_bits[15519:15488];
                // 10'h1e5 :  sha3_din <= random_bits[15551:15520];
                // 10'h1e6 :  sha3_din <= random_bits[15583:15552];
                // 10'h1e7 :  sha3_din <= random_bits[15615:15584];
                // 10'h1e8 :  sha3_din <= random_bits[15647:15616];
                // 10'h1e9 :  sha3_din <= random_bits[15679:15648];
                // 10'h1ea :  sha3_din <= random_bits[15711:15680];
                // 10'h1eb :  sha3_din <= random_bits[15743:15712];
                // 10'h1ec :  sha3_din <= random_bits[15775:15744];
                // 10'h1ed :  sha3_din <= random_bits[15807:15776];
                // 10'h1ee :  sha3_din <= random_bits[15839:15808];
                // 10'h1ef :  sha3_din <= random_bits[15871:15840];
                // 10'h1f0 :  sha3_din <= random_bits[15903:15872];
                // 10'h1f1 :  sha3_din <= random_bits[15935:15904];
                // 10'h1f2 :  sha3_din <= random_bits[15967:15936];
                // 10'h1f3 :  sha3_din <= random_bits[15999:15968];
                // 10'h1f4 :  sha3_din <= random_bits[16031:16000];
                // 10'h1f5 :  sha3_din <= random_bits[16063:16032];
                // 10'h1f6 :  sha3_din <= random_bits[16095:16064];
                // 10'h1f7 :  sha3_din <= random_bits[16127:16096];
                // 10'h1f8 :  sha3_din <= random_bits[16159:16128];
                // 10'h1f9 :  sha3_din <= random_bits[16191:16160];
                // 10'h1fa :  sha3_din <= random_bits[16223:16192];
                // 10'h1fb :  sha3_din <= random_bits[16255:16224];
                // 10'h1fc :  sha3_din <= random_bits[16287:16256];
                // 10'h1fd :  sha3_din <= random_bits[16319:16288];
                // 10'h1fe :  sha3_din <= random_bits[16351:16320];
                // 10'h1ff :  sha3_din <= random_bits[16383:16352];
                // 10'h200 :  sha3_din <= random_bits[16415:16384];
                // 10'h201 :  sha3_din <= random_bits[16447:16416];
                // 10'h202 :  sha3_din <= random_bits[16479:16448];
                // 10'h203 :  sha3_din <= random_bits[16511:16480];
                // 10'h204 :  sha3_din <= random_bits[16543:16512];
                // 10'h205 :  sha3_din <= random_bits[16575:16544];
                // 10'h206 :  sha3_din <= random_bits[16607:16576];
                // 10'h207 :  sha3_din <= random_bits[16639:16608];
                // 10'h208 :  sha3_din <= random_bits[16671:16640];
                // 10'h209 :  sha3_din <= random_bits[16703:16672];
                // 10'h20a :  sha3_din <= random_bits[16735:16704];
                // 10'h20b :  sha3_din <= random_bits[16767:16736];
                // 10'h20c :  sha3_din <= random_bits[16799:16768];
                // 10'h20d :  sha3_din <= random_bits[16831:16800];
                // 10'h20e :  sha3_din <= random_bits[16863:16832];
                // 10'h20f :  sha3_din <= random_bits[16895:16864];
                // 10'h210 :  sha3_din <= random_bits[16927:16896];
                // 10'h211 :  sha3_din <= random_bits[16959:16928];
                // 10'h212 :  sha3_din <= random_bits[16991:16960];
                // 10'h213 :  sha3_din <= random_bits[17023:16992];
                // 10'h214 :  sha3_din <= random_bits[17055:17024];
                // 10'h215 :  sha3_din <= random_bits[17087:17056];
                // 10'h216 :  sha3_din <= random_bits[17119:17088];
                // 10'h217 :  sha3_din <= random_bits[17151:17120];
                // 10'h218 :  sha3_din <= random_bits[17183:17152];
                // 10'h219 :  sha3_din <= random_bits[17215:17184];
                // 10'h21a :  sha3_din <= random_bits[17247:17216];
                // 10'h21b :  sha3_din <= random_bits[17279:17248];
                // 10'h21c :  sha3_din <= random_bits[17311:17280];
                // 10'h21d :  sha3_din <= random_bits[17343:17312];
                // 10'h21e :  sha3_din <= random_bits[17375:17344];
                // 10'h21f :  sha3_din <= random_bits[17407:17376];
                // 10'h220 :  sha3_din <= random_bits[17439:17408];
                // 10'h221 :  sha3_din <= random_bits[17471:17440];
                // 10'h222 :  sha3_din <= random_bits[17503:17472];
                // 10'h223 :  sha3_din <= random_bits[17535:17504];
                // 10'h224 :  sha3_din <= random_bits[17567:17536];
                // 10'h225 :  sha3_din <= random_bits[17599:17568];
                // 10'h226 :  sha3_din <= random_bits[17631:17600];
                // 10'h227 :  sha3_din <= random_bits[17663:17632];
                // 10'h228 :  sha3_din <= random_bits[17695:17664];
                // 10'h229 :  sha3_din <= random_bits[17727:17696];
                // 10'h22a :  sha3_din <= random_bits[17759:17728];
                // 10'h22b :  sha3_din <= random_bits[17791:17760];
                // 10'h22c :  sha3_din <= random_bits[17823:17792];
                // 10'h22d :  sha3_din <= random_bits[17855:17824];
                // 10'h22e :  sha3_din <= random_bits[17887:17856];
                // 10'h22f :  sha3_din <= random_bits[17919:17888];
                // 10'h230 :  sha3_din <= random_bits[17951:17920];
                // 10'h231 :  sha3_din <= random_bits[17983:17952];
                // 10'h232 :  sha3_din <= random_bits[18015:17984];
                // 10'h233 :  sha3_din <= random_bits[18047:18016];
                // 10'h234 :  sha3_din <= random_bits[18079:18048];
                // 10'h235 :  sha3_din <= random_bits[18111:18080];
                // 10'h236 :  sha3_din <= random_bits[18143:18112];
                // 10'h237 :  sha3_din <= random_bits[18175:18144];
                // 10'h238 :  sha3_din <= random_bits[18207:18176];
                // 10'h239 :  sha3_din <= random_bits[18239:18208];
                // 10'h23a :  sha3_din <= random_bits[18271:18240];
                // 10'h23b :  sha3_din <= random_bits[18303:18272];
                // 10'h23c :  sha3_din <= random_bits[18335:18304];
                // 10'h23d :  sha3_din <= random_bits[18367:18336];
                // 10'h23e :  sha3_din <= random_bits[18399:18368];
                // 10'h23f :  sha3_din <= random_bits[18431:18400];
                // 10'h240 :  sha3_din <= random_bits[18463:18432];
                // 10'h241 :  sha3_din <= random_bits[18495:18464];
                // 10'h242 :  sha3_din <= random_bits[18527:18496];
                // 10'h243 :  sha3_din <= random_bits[18559:18528];
                // 10'h244 :  sha3_din <= random_bits[18591:18560];
                // 10'h245 :  sha3_din <= random_bits[18623:18592];
                // 10'h246 :  sha3_din <= random_bits[18655:18624];
                // 10'h247 :  sha3_din <= random_bits[18687:18656];
                // 10'h248 :  sha3_din <= random_bits[18719:18688];
                // 10'h249 :  sha3_din <= random_bits[18751:18720];
                // 10'h24a :  sha3_din <= random_bits[18783:18752];
                // 10'h24b :  sha3_din <= random_bits[18815:18784];
                // 10'h24c :  sha3_din <= random_bits[18847:18816];
                // 10'h24d :  sha3_din <= random_bits[18879:18848];
                // 10'h24e :  sha3_din <= random_bits[18911:18880];
                // 10'h24f :  sha3_din <= random_bits[18943:18912];
                // 10'h250 :  sha3_din <= random_bits[18975:18944];
                // 10'h251 :  sha3_din <= random_bits[19007:18976];
                // 10'h252 :  sha3_din <= random_bits[19039:19008];
                // 10'h253 :  sha3_din <= random_bits[19071:19040];
                // 10'h254 :  sha3_din <= random_bits[19103:19072];
                // 10'h255 :  sha3_din <= random_bits[19135:19104];
                // 10'h256 :  sha3_din <= random_bits[19167:19136];
                // 10'h257 :  sha3_din <= random_bits[19199:19168];
                // 10'h258 :  sha3_din <= random_bits[19231:19200];
                // 10'h259 :  sha3_din <= random_bits[19263:19232];
                // 10'h25a :  sha3_din <= random_bits[19295:19264];
                // 10'h25b :  sha3_din <= random_bits[19327:19296];
                // 10'h25c :  sha3_din <= random_bits[19359:19328];
                // 10'h25d :  sha3_din <= random_bits[19391:19360];
                // 10'h25e :  sha3_din <= random_bits[19423:19392];
                // 10'h25f :  sha3_din <= random_bits[19455:19424];
                // 10'h260 :  sha3_din <= random_bits[19487:19456];
                // 10'h261 :  sha3_din <= random_bits[19519:19488];
                // 10'h262 :  sha3_din <= random_bits[19551:19520];
                // 10'h263 :  sha3_din <= random_bits[19583:19552];
                // 10'h264 :  sha3_din <= random_bits[19615:19584];
                // 10'h265 :  sha3_din <= random_bits[19647:19616];
                // 10'h266 :  sha3_din <= random_bits[19679:19648];
                // 10'h267 :  sha3_din <= random_bits[19711:19680];
                // 10'h268 :  sha3_din <= random_bits[19743:19712];
                // 10'h269 :  sha3_din <= random_bits[19775:19744];
                // 10'h26a :  sha3_din <= random_bits[19807:19776];
                // 10'h26b :  sha3_din <= random_bits[19839:19808];
                // 10'h26c :  sha3_din <= random_bits[19871:19840];
                // 10'h26d :  sha3_din <= random_bits[19903:19872];
                // 10'h26e :  sha3_din <= random_bits[19935:19904];
                // 10'h26f :  sha3_din <= random_bits[19967:19936];
                // 10'h270 :  sha3_din <= random_bits[19999:19968];
                // 10'h271 :  sha3_din <= random_bits[20031:20000];
                // 10'h272 :  sha3_din <= random_bits[20063:20032];
                // 10'h273 :  sha3_din <= random_bits[20095:20064];
                // 10'h274 :  sha3_din <= random_bits[20127:20096];
                // 10'h275 :  sha3_din <= random_bits[20159:20128];
                // 10'h276 :  sha3_din <= random_bits[20191:20160];
                // 10'h277 :  sha3_din <= random_bits[20223:20192];
                // 10'h278 :  sha3_din <= random_bits[20255:20224];
                // 10'h279 :  sha3_din <= random_bits[20287:20256];
                // 10'h27a :  sha3_din <= random_bits[20319:20288];
                // 10'h27b :  sha3_din <= random_bits[20351:20320];
                // 10'h27c :  sha3_din <= random_bits[20383:20352];
                // 10'h27d :  sha3_din <= random_bits[20415:20384];
                // 10'h27e :  sha3_din <= random_bits[20447:20416];
                // 10'h27f :  sha3_din <= random_bits[20479:20448];
                // 10'h280 :  sha3_din <= random_bits[20511:20480];
                // 10'h281 :  sha3_din <= random_bits[20543:20512];
                // 10'h282 :  sha3_din <= random_bits[20575:20544];
                // 10'h283 :  sha3_din <= random_bits[20607:20576];
                // 10'h284 :  sha3_din <= random_bits[20639:20608];
                // 10'h285 :  sha3_din <= random_bits[20671:20640];
                // 10'h286 :  sha3_din <= random_bits[20703:20672];
                // 10'h287 :  sha3_din <= random_bits[20735:20704];
                // 10'h288 :  sha3_din <= random_bits[20767:20736];
                // 10'h289 :  sha3_din <= random_bits[20799:20768];
                // 10'h28a :  sha3_din <= random_bits[20831:20800];
                // 10'h28b :  sha3_din <= random_bits[20863:20832];
                // 10'h28c :  sha3_din <= random_bits[20895:20864];
                // 10'h28d :  sha3_din <= random_bits[20927:20896];
                // 10'h28e :  sha3_din <= random_bits[20959:20928];
                // 10'h28f :  sha3_din <= random_bits[20991:20960];
                // 10'h290 :  sha3_din <= random_bits[21023:20992];
                // 10'h291 :  sha3_din <= random_bits[21055:21024];
                // 10'h292 :  sha3_din <= random_bits[21087:21056];
                // 10'h293 :  sha3_din <= random_bits[21119:21088];
                // 10'h294 :  sha3_din <= random_bits[21151:21120];
                // 10'h295 :  sha3_din <= random_bits[21183:21152];
                // 10'h296 :  sha3_din <= random_bits[21215:21184];
                // 10'h297 :  sha3_din <= random_bits[21247:21216];
                // 10'h298 :  sha3_din <= random_bits[21279:21248];
                // 10'h299 :  sha3_din <= random_bits[21311:21280];
                // 10'h29a :  sha3_din <= random_bits[21343:21312];
                // 10'h29b :  sha3_din <= random_bits[21375:21344];
                // 10'h29c :  sha3_din <= random_bits[21407:21376];
                // 10'h29d :  sha3_din <= random_bits[21439:21408];
                // 10'h29e :  sha3_din <= random_bits[21471:21440];
                // 10'h29f :  sha3_din <= random_bits[21503:21472];
                // 10'h2a0 :  sha3_din <= random_bits[21535:21504];
                // 10'h2a1 :  sha3_din <= random_bits[21567:21536];
                // 10'h2a2 :  sha3_din <= random_bits[21599:21568];
                // 10'h2a3 :  sha3_din <= random_bits[21631:21600];
                // 10'h2a4 :  sha3_din <= random_bits[21663:21632];
                // 10'h2a5 :  sha3_din <= random_bits[21695:21664];
                // 10'h2a6 :  sha3_din <= random_bits[21727:21696];
                // 10'h2a7 :  sha3_din <= random_bits[21759:21728];
                // 10'h2a8 :  sha3_din <= random_bits[21791:21760];
                // 10'h2a9 :  sha3_din <= random_bits[21823:21792];
                // 10'h2aa :  sha3_din <= random_bits[21855:21824];
                // 10'h2ab :  sha3_din <= random_bits[21887:21856];
                // 10'h2ac :  sha3_din <= random_bits[21919:21888];
                // 10'h2ad :  sha3_din <= random_bits[21951:21920];
                // 10'h2ae :  sha3_din <= random_bits[21983:21952];
                // 10'h2af :  sha3_din <= random_bits[22015:21984];
                // 10'h2b0 :  sha3_din <= random_bits[22047:22016];
                // 10'h2b1 :  sha3_din <= random_bits[22079:22048];
                // 10'h2b2 :  sha3_din <= random_bits[22111:22080];
                // 10'h2b3 :  sha3_din <= random_bits[22143:22112];
                // 10'h2b4 :  sha3_din <= random_bits[22175:22144];
                // 10'h2b5 :  sha3_din <= random_bits[22207:22176];
                // 10'h2b6 :  sha3_din <= random_bits[22239:22208];
                // 10'h2b7 :  sha3_din <= random_bits[22271:22240];
                // 10'h2b8 :  sha3_din <= random_bits[22303:22272];
                // 10'h2b9 :  sha3_din <= random_bits[22335:22304];
                // 10'h2ba :  sha3_din <= random_bits[22367:22336];
                // 10'h2bb :  sha3_din <= random_bits[22399:22368];
                // 10'h2bc :  sha3_din <= random_bits[22431:22400];
                // 10'h2bd :  sha3_din <= random_bits[22463:22432];
                // 10'h2be :  sha3_din <= random_bits[22495:22464];
                // 10'h2bf :  sha3_din <= random_bits[22527:22496];
                // 10'h2c0 :  sha3_din <= random_bits[22559:22528];
                // 10'h2c1 :  sha3_din <= random_bits[22591:22560];
                // 10'h2c2 :  sha3_din <= random_bits[22623:22592];
                // 10'h2c3 :  sha3_din <= random_bits[22655:22624];
                // 10'h2c4 :  sha3_din <= random_bits[22687:22656];
                // 10'h2c5 :  sha3_din <= random_bits[22719:22688];
                // 10'h2c6 :  sha3_din <= random_bits[22751:22720];
                // 10'h2c7 :  sha3_din <= random_bits[22783:22752];
                // 10'h2c8 :  sha3_din <= random_bits[22815:22784];
                // 10'h2c9 :  sha3_din <= random_bits[22847:22816];
                // 10'h2ca :  sha3_din <= random_bits[22879:22848];
                // 10'h2cb :  sha3_din <= random_bits[22911:22880];
                // 10'h2cc :  sha3_din <= random_bits[22943:22912];
                // 10'h2cd :  sha3_din <= random_bits[22975:22944];
                // 10'h2ce :  sha3_din <= random_bits[23007:22976];
                // 10'h2cf :  sha3_din <= random_bits[23039:23008];
                // 10'h2d0 :  sha3_din <= random_bits[23071:23040];
                // 10'h2d1 :  sha3_din <= random_bits[23103:23072];
                // 10'h2d2 :  sha3_din <= random_bits[23135:23104];
                // 10'h2d3 :  sha3_din <= random_bits[23167:23136];
                // 10'h2d4 :  sha3_din <= random_bits[23199:23168];
                // 10'h2d5 :  sha3_din <= random_bits[23231:23200];
                // 10'h2d6 :  sha3_din <= random_bits[23263:23232];
                // 10'h2d7 :  sha3_din <= random_bits[23295:23264];
                // 10'h2d8 :  sha3_din <= random_bits[23327:23296];
                // 10'h2d9 :  sha3_din <= random_bits[23359:23328];
                // 10'h2da :  sha3_din <= random_bits[23391:23360];
                // 10'h2db :  sha3_din <= random_bits[23423:23392];
                // 10'h2dc :  sha3_din <= random_bits[23455:23424];
                // 10'h2dd :  sha3_din <= random_bits[23487:23456];
                // 10'h2de :  sha3_din <= random_bits[23519:23488];
                // 10'h2df :  sha3_din <= random_bits[23551:23520];
                // 10'h2e0 :  sha3_din <= random_bits[23583:23552];
                // 10'h2e1 :  sha3_din <= random_bits[23615:23584];
                // 10'h2e2 :  sha3_din <= random_bits[23647:23616];
                // 10'h2e3 :  sha3_din <= random_bits[23679:23648];
                // 10'h2e4 :  sha3_din <= random_bits[23711:23680];
                // 10'h2e5 :  sha3_din <= random_bits[23743:23712];
                // 10'h2e6 :  sha3_din <= random_bits[23775:23744];
                // 10'h2e7 :  sha3_din <= random_bits[23807:23776];
                // 10'h2e8 :  sha3_din <= random_bits[23839:23808];
                // 10'h2e9 :  sha3_din <= random_bits[23871:23840];
                // 10'h2ea :  sha3_din <= random_bits[23903:23872];
                // 10'h2eb :  sha3_din <= random_bits[23935:23904];
                // 10'h2ec :  sha3_din <= random_bits[23967:23936];
                // 10'h2ed :  sha3_din <= random_bits[23999:23968];
                // 10'h2ee :  sha3_din <= random_bits[24031:24000];
                // 10'h2ef :  sha3_din <= random_bits[24063:24032];
                // 10'h2f0 :  sha3_din <= random_bits[24095:24064];
                // 10'h2f1 :  sha3_din <= random_bits[24127:24096];
                // 10'h2f2 :  sha3_din <= random_bits[24159:24128];
                // 10'h2f3 :  sha3_din <= random_bits[24191:24160];
                // 10'h2f4 :  sha3_din <= random_bits[24223:24192];
                // 10'h2f5 :  sha3_din <= random_bits[24255:24224];
                // 10'h2f6 :  sha3_din <= random_bits[24287:24256];
                // 10'h2f7 :  sha3_din <= random_bits[24319:24288];
                // 10'h2f8 :  sha3_din <= random_bits[24351:24320];
                // 10'h2f9 :  sha3_din <= random_bits[24383:24352];
                // 10'h2fa :  sha3_din <= random_bits[24415:24384];
                // 10'h2fb :  sha3_din <= random_bits[24447:24416];
                // 10'h2fc :  sha3_din <= random_bits[24479:24448];
                // 10'h2fd :  sha3_din <= random_bits[24511:24480];
                // 10'h2fe :  sha3_din <= random_bits[24543:24512];
                // 10'h2ff :  sha3_din <= random_bits[24575:24544];
                // 10'h300 :  sha3_din <= random_bits[24607:24576];
                // 10'h301 :  sha3_din <= random_bits[24639:24608];
                // 10'h302 :  sha3_din <= random_bits[24671:24640];
                // 10'h303 :  sha3_din <= random_bits[24703:24672];
                // 10'h304 :  sha3_din <= random_bits[24735:24704];
                // 10'h305 :  sha3_din <= random_bits[24767:24736];
                // 10'h306 :  sha3_din <= random_bits[24799:24768];
                // 10'h307 :  sha3_din <= random_bits[24831:24800];
                // 10'h308 :  sha3_din <= random_bits[24863:24832];
                // 10'h309 :  sha3_din <= random_bits[24895:24864];
                // 10'h30a :  sha3_din <= random_bits[24927:24896];
                // 10'h30b :  sha3_din <= random_bits[24959:24928];
                // 10'h30c :  sha3_din <= random_bits[24991:24960];
                // 10'h30d :  sha3_din <= random_bits[25023:24992];
                // 10'h30e :  sha3_din <= random_bits[25055:25024];
                // 10'h30f :  sha3_din <= random_bits[25087:25056];
                // 10'h310 :  sha3_din <= random_bits[25119:25088];
                // 10'h311 :  sha3_din <= random_bits[25151:25120];
                // 10'h312 :  sha3_din <= random_bits[25183:25152];
                // 10'h313 :  sha3_din <= random_bits[25215:25184];
                // 10'h314 :  sha3_din <= random_bits[25247:25216];
                // 10'h315 :  sha3_din <= random_bits[25279:25248];
                // 10'h316 :  sha3_din <= random_bits[25311:25280];
                // 10'h317 :  sha3_din <= random_bits[25343:25312];
                // 10'h318 :  sha3_din <= random_bits[25375:25344];
                // 10'h319 :  sha3_din <= random_bits[25407:25376];
                // 10'h31a :  sha3_din <= random_bits[25439:25408];
                // 10'h31b :  sha3_din <= random_bits[25471:25440];
                // 10'h31c :  sha3_din <= random_bits[25503:25472];
                // 10'h31d :  sha3_din <= random_bits[25535:25504];
                // 10'h31e :  sha3_din <= random_bits[25567:25536];
                // 10'h31f :  sha3_din <= random_bits[25599:25568];
                // 10'h320 :  sha3_din <= random_bits[25631:25600];
                // 10'h321 :  sha3_din <= random_bits[25663:25632];
                // 10'h322 :  sha3_din <= random_bits[25695:25664];
                // 10'h323 :  sha3_din <= random_bits[25727:25696];
                // 10'h324 :  sha3_din <= random_bits[25759:25728];
                // 10'h325 :  sha3_din <= random_bits[25791:25760];
                // 10'h326 :  sha3_din <= random_bits[25823:25792];
                // 10'h327 :  sha3_din <= random_bits[25855:25824];
                // 10'h328 :  sha3_din <= random_bits[25887:25856];
                // 10'h329 :  sha3_din <= random_bits[25919:25888];
                // 10'h32a :  sha3_din <= random_bits[25951:25920];
                // 10'h32b :  sha3_din <= random_bits[25983:25952];
                // 10'h32c :  sha3_din <= random_bits[26015:25984];
                // 10'h32d :  sha3_din <= random_bits[26047:26016];
                // 10'h32e :  sha3_din <= random_bits[26079:26048];
                // 10'h32f :  sha3_din <= random_bits[26111:26080];
                // 10'h330 :  sha3_din <= random_bits[26143:26112];
                // 10'h331 :  sha3_din <= random_bits[26175:26144];
                // 10'h332 :  sha3_din <= random_bits[26207:26176];
                // 10'h333 :  sha3_din <= random_bits[26239:26208];
                // 10'h334 :  sha3_din <= random_bits[26271:26240];
                // 10'h335 :  sha3_din <= random_bits[26303:26272];
                // 10'h336 :  sha3_din <= random_bits[26335:26304];
                // 10'h337 :  sha3_din <= random_bits[26367:26336];
                // 10'h338 :  sha3_din <= random_bits[26399:26368];
                // 10'h339 :  sha3_din <= random_bits[26431:26400];
                // 10'h33a :  sha3_din <= random_bits[26463:26432];
                // 10'h33b :  sha3_din <= random_bits[26495:26464];
                // 10'h33c :  sha3_din <= random_bits[26527:26496];
                // 10'h33d :  sha3_din <= random_bits[26559:26528];
                // 10'h33e :  sha3_din <= random_bits[26591:26560];
                // 10'h33f :  sha3_din <= random_bits[26623:26592];
                // 10'h340 :  sha3_din <= random_bits[26655:26624];
                // 10'h341 :  sha3_din <= random_bits[26687:26656];
                // 10'h342 :  sha3_din <= random_bits[26719:26688];
                // 10'h343 :  sha3_din <= random_bits[26751:26720];
                // 10'h344 :  sha3_din <= random_bits[26783:26752];
                // 10'h345 :  sha3_din <= random_bits[26815:26784];
                // 10'h346 :  sha3_din <= random_bits[26847:26816];
                // 10'h347 :  sha3_din <= random_bits[26879:26848];
                // 10'h348 :  sha3_din <= random_bits[26911:26880];
                // 10'h349 :  sha3_din <= random_bits[26943:26912];
                // 10'h34a :  sha3_din <= random_bits[26975:26944];
                // 10'h34b :  sha3_din <= random_bits[27007:26976];
                // 10'h34c :  sha3_din <= random_bits[27039:27008];
                // 10'h34d :  sha3_din <= random_bits[27071:27040];
                // 10'h34e :  sha3_din <= random_bits[27103:27072];
                // 10'h34f :  sha3_din <= random_bits[27135:27104];
                // 10'h350 :  sha3_din <= random_bits[27167:27136];
                // 10'h351 :  sha3_din <= random_bits[27199:27168];
                // 10'h352 :  sha3_din <= random_bits[27231:27200];
                // 10'h353 :  sha3_din <= random_bits[27263:27232];
                // 10'h354 :  sha3_din <= random_bits[27295:27264];
                // 10'h355 :  sha3_din <= random_bits[27327:27296];
                // 10'h356 :  sha3_din <= random_bits[27359:27328];
                // 10'h357 :  sha3_din <= random_bits[27391:27360];
                // 10'h358 :  sha3_din <= random_bits[27423:27392];
                // 10'h359 :  sha3_din <= random_bits[27455:27424];
                // 10'h35a :  sha3_din <= random_bits[27487:27456];
                // 10'h35b :  sha3_din <= random_bits[27519:27488];
                // 10'h35c :  sha3_din <= random_bits[27551:27520];
                // 10'h35d :  sha3_din <= random_bits[27583:27552];
                // 10'h35e :  sha3_din <= random_bits[27615:27584];
                // 10'h35f :  sha3_din <= random_bits[27647:27616];
                // 10'h360 :  sha3_din <= random_bits[27679:27648];
                // 10'h361 :  sha3_din <= random_bits[27711:27680];
                // 10'h362 :  sha3_din <= random_bits[27743:27712];
                // 10'h363 :  sha3_din <= random_bits[27775:27744];
                // 10'h364 :  sha3_din <= random_bits[27807:27776];
                // 10'h365 :  sha3_din <= random_bits[27839:27808];
                // 10'h366 :  sha3_din <= random_bits[27871:27840];
                // 10'h367 :  sha3_din <= random_bits[27903:27872];
                // 10'h368 :  sha3_din <= random_bits[27935:27904];
                // 10'h369 :  sha3_din <= random_bits[27967:27936];
                // 10'h36a :  sha3_din <= random_bits[27999:27968];
                // 10'h36b :  sha3_din <= random_bits[28031:28000];
                // 10'h36c :  sha3_din <= random_bits[28063:28032];
                // 10'h36d :  sha3_din <= random_bits[28095:28064];
                // 10'h36e :  sha3_din <= random_bits[28127:28096];
                // 10'h36f :  sha3_din <= random_bits[28159:28128];
                // 10'h370 :  sha3_din <= random_bits[28191:28160];
                // 10'h371 :  sha3_din <= random_bits[28223:28192];
                // 10'h372 :  sha3_din <= random_bits[28255:28224];
                // 10'h373 :  sha3_din <= random_bits[28287:28256];
                // 10'h374 :  sha3_din <= random_bits[28319:28288];
                // 10'h375 :  sha3_din <= random_bits[28351:28320];
                // 10'h376 :  sha3_din <= random_bits[28383:28352];
                // 10'h377 :  sha3_din <= random_bits[28415:28384];
                // 10'h378 :  sha3_din <= random_bits[28447:28416];
                // 10'h379 :  sha3_din <= random_bits[28479:28448];
                // 10'h37a :  sha3_din <= random_bits[28511:28480];
                // 10'h37b :  sha3_din <= random_bits[28543:28512];
                // 10'h37c :  sha3_din <= random_bits[28575:28544];
                // 10'h37d :  sha3_din <= random_bits[28607:28576];
                // 10'h37e :  sha3_din <= random_bits[28639:28608];
                // 10'h37f :  sha3_din <= random_bits[28671:28640];
                // 10'h380 :  sha3_din <= random_bits[28703:28672];
                // 10'h381 :  sha3_din <= random_bits[28735:28704];
                // 10'h382 :  sha3_din <= random_bits[28767:28736];
                // 10'h383 :  sha3_din <= random_bits[28799:28768];
                // 10'h384 :  sha3_din <= random_bits[28831:28800];
                // 10'h385 :  sha3_din <= random_bits[28863:28832];
                // 10'h386 :  sha3_din <= random_bits[28895:28864];
                // 10'h387 :  sha3_din <= random_bits[28927:28896];
                // 10'h388 :  sha3_din <= random_bits[28959:28928];
                // 10'h389 :  sha3_din <= random_bits[28991:28960];
                // 10'h38a :  sha3_din <= random_bits[29023:28992];
                // 10'h38b :  sha3_din <= random_bits[29055:29024];
                // 10'h38c :  sha3_din <= random_bits[29087:29056];
                // 10'h38d :  sha3_din <= random_bits[29119:29088];
                // 10'h38e :  sha3_din <= random_bits[29151:29120];
                // 10'h38f :  sha3_din <= random_bits[29183:29152];
                // 10'h390 :  sha3_din <= random_bits[29215:29184];
                // 10'h391 :  sha3_din <= random_bits[29247:29216];
                // 10'h392 :  sha3_din <= random_bits[29279:29248];
                // 10'h393 :  sha3_din <= random_bits[29311:29280];
                // 10'h394 :  sha3_din <= random_bits[29343:29312];
                // 10'h395 :  sha3_din <= random_bits[29375:29344];
                // 10'h396 :  sha3_din <= random_bits[29407:29376];
                // 10'h397 :  sha3_din <= random_bits[29439:29408];
                // 10'h398 :  sha3_din <= random_bits[29471:29440];
                // 10'h399 :  sha3_din <= random_bits[29503:29472];
                // 10'h39a :  sha3_din <= random_bits[29535:29504];
                // 10'h39b :  sha3_din <= random_bits[29567:29536];
                // 10'h39c :  sha3_din <= random_bits[29599:29568];
                // 10'h39d :  sha3_din <= random_bits[29631:29600];
                // 10'h39e :  sha3_din <= random_bits[29663:29632];
                // 10'h39f :  sha3_din <= random_bits[29695:29664];
                // 10'h3a0 :  sha3_din <= random_bits[29727:29696];
                // 10'h3a1 :  sha3_din <= random_bits[29759:29728];
                // 10'h3a2 :  sha3_din <= random_bits[29791:29760];
                // 10'h3a3 :  sha3_din <= random_bits[29823:29792];
                // 10'h3a4 :  sha3_din <= random_bits[29855:29824];
                // 10'h3a5 :  sha3_din <= random_bits[29887:29856];
                // 10'h3a6 :  sha3_din <= random_bits[29919:29888];
                // 10'h3a7 :  sha3_din <= random_bits[29951:29920];
                // 10'h3a8 :  sha3_din <= random_bits[29983:29952];
                // 10'h3a9 :  sha3_din <= random_bits[30015:29984];
                // 10'h3aa :  sha3_din <= random_bits[30047:30016];
                // 10'h3ab :  sha3_din <= random_bits[30079:30048];
                // 10'h3ac :  sha3_din <= random_bits[30111:30080];
                // 10'h3ad :  sha3_din <= random_bits[30143:30112];
                // 10'h3ae :  sha3_din <= random_bits[30175:30144];
                // 10'h3af :  sha3_din <= random_bits[30207:30176];
                // 10'h3b0 :  sha3_din <= random_bits[30239:30208];
                // 10'h3b1 :  sha3_din <= random_bits[30271:30240];
                // 10'h3b2 :  sha3_din <= random_bits[30303:30272];
                // 10'h3b3 :  sha3_din <= random_bits[30335:30304];
                // 10'h3b4 :  sha3_din <= random_bits[30367:30336];
                // 10'h3b5 :  sha3_din <= random_bits[30399:30368];
                // 10'h3b6 :  sha3_din <= random_bits[30431:30400];
                // 10'h3b7 :  sha3_din <= random_bits[30463:30432];
                // 10'h3b8 :  sha3_din <= random_bits[30495:30464];
                // 10'h3b9 :  sha3_din <= random_bits[30527:30496];
                // 10'h3ba :  sha3_din <= random_bits[30559:30528];
                // 10'h3bb :  sha3_din <= random_bits[30591:30560];
                // 10'h3bc :  sha3_din <= random_bits[30623:30592];
                // 10'h3bd :  sha3_din <= random_bits[30655:30624];
                // 10'h3be :  sha3_din <= random_bits[30687:30656];
                // 10'h3bf :  sha3_din <= random_bits[30719:30688];
                // 10'h3c0 :  sha3_din <= random_bits[30751:30720];
                // 10'h3c1 :  sha3_din <= random_bits[30783:30752];
                // 10'h3c2 :  sha3_din <= random_bits[30815:30784];
                // 10'h3c3 :  sha3_din <= random_bits[30847:30816];
                // 10'h3c4 :  sha3_din <= random_bits[30879:30848];
                // 10'h3c5 :  sha3_din <= random_bits[30911:30880];
                // 10'h3c6 :  sha3_din <= random_bits[30943:30912];
                // 10'h3c7 :  sha3_din <= random_bits[30975:30944];
                // 10'h3c8 :  sha3_din <= random_bits[31007:30976];
                // 10'h3c9 :  sha3_din <= random_bits[31039:31008];
                // 10'h3ca :  sha3_din <= random_bits[31071:31040];
                // 10'h3cb :  sha3_din <= random_bits[31103:31072];
                // 10'h3cc :  sha3_din <= random_bits[31135:31104];
                // 10'h3cd :  sha3_din <= random_bits[31167:31136];
                // 10'h3ce :  sha3_din <= random_bits[31199:31168];
                // 10'h3cf :  sha3_din <= random_bits[31231:31200];
                // 10'h3d0 :  sha3_din <= random_bits[31263:31232];
                // 10'h3d1 :  sha3_din <= random_bits[31295:31264];
                // 10'h3d2 :  sha3_din <= random_bits[31327:31296];
                // 10'h3d3 :  sha3_din <= random_bits[31359:31328];
                // 10'h3d4 :  sha3_din <= random_bits[31391:31360];
                // 10'h3d5 :  sha3_din <= random_bits[31423:31392];
                // 10'h3d6 :  sha3_din <= random_bits[31455:31424];
                // 10'h3d7 :  sha3_din <= random_bits[31487:31456];
                // 10'h3d8 :  sha3_din <= random_bits[31519:31488];
                // 10'h3d9 :  sha3_din <= random_bits[31551:31520];
                // 10'h3da :  sha3_din <= random_bits[31583:31552];
                // 10'h3db :  sha3_din <= random_bits[31615:31584];
                // 10'h3dc :  sha3_din <= random_bits[31647:31616];
                // 10'h3dd :  sha3_din <= random_bits[31679:31648];
                // 10'h3de :  sha3_din <= random_bits[31711:31680];
                // 10'h3df :  sha3_din <= random_bits[31743:31712];
                // 10'h3e0 :  sha3_din <= random_bits[31775:31744];
                // 10'h3e1 :  sha3_din <= random_bits[31807:31776];
                // 10'h3e2 :  sha3_din <= random_bits[31839:31808];
                // 10'h3e3 :  sha3_din <= random_bits[31871:31840];
                // 10'h3e4 :  sha3_din <= random_bits[31903:31872];
                // 10'h3e5 :  sha3_din <= random_bits[31935:31904];
                // 10'h3e6 :  sha3_din <= random_bits[31967:31936];
                // 10'h3e7 :  sha3_din <= random_bits[31999:31968];
                // 10'h3e8 :  sha3_din <= random_bits[32031:32000];
                // 10'h3e9 :  sha3_din <= random_bits[32063:32032];
                // 10'h3ea :  sha3_din <= random_bits[32095:32064];
                // 10'h3eb :  sha3_din <= random_bits[32127:32096];
                // 10'h3ec :  sha3_din <= random_bits[32159:32128];
                // 10'h3ed :  sha3_din <= random_bits[32191:32160];
                // 10'h3ee :  sha3_din <= random_bits[32223:32192];
                // 10'h3ef :  sha3_din <= random_bits[32255:32224];
                // 10'h3f0 :  sha3_din <= random_bits[32287:32256];
                // 10'h3f1 :  sha3_din <= random_bits[32319:32288];
                // 10'h3f2 :  sha3_din <= random_bits[32351:32320];
                // 10'h3f3 :  sha3_din <= random_bits[32383:32352];
                // 10'h3f4 :  sha3_din <= random_bits[32415:32384];
                // 10'h3f5 :  sha3_din <= random_bits[32447:32416];
                // 10'h3f6 :  sha3_din <= random_bits[32479:32448];
                // 10'h3f7 :  sha3_din <= random_bits[32511:32480];
                // 10'h3f8 :  sha3_din <= random_bits[32543:32512];
                // 10'h3f9 :  sha3_din <= random_bits[32575:32544];
                // 10'h3fa :  sha3_din <= random_bits[32607:32576];
                // 10'h3fb :  sha3_din <= random_bits[32639:32608];
                // 10'h3fc :  sha3_din <= random_bits[32671:32640];
                // 10'h3fd :  sha3_din <= random_bits[32703:32672];
                // 10'h3fe :  sha3_din <= random_bits[32735:32704];
                // 10'h3ff :  sha3_din <= random_bits[32767:32736];
                default :  sha3_din <= random_bits[31:0];
            endcase
            writed_words_counter <= writed_words_counter + 1;
            sha3_we  <= 1;
            //sha3_cs <= 1;
            //sha3_cs <= 1;
            if(writed_words_counter  == NUMBER_OF_WORDS_SHA3INIT)
            begin
                state <= writed_to_sha ;
                writed_words_counter  <= 0; 
            end
         end
         
         writed_to_sha: begin//dane zapisane ////4
            sha3_we <= 0;//opuszczenie flag zapisania do wewnętrznego rejestru
            sha3_address <= 0;
            sha3_din  <= 0;
            //TODO! w zależności, czy blok pierwszy czy kolejny zmienić
            sha3_init <= 1;
            state <= generating_hash;
            
//            if(writed_words_counter == 8'hFF)
//            begin
//                state <= final_hash_generation;
//            end
//            else if(writed_words_counter_mod16  == 8'h00)
//            begin
//                state <= generating_hash;
//            end
//            else
//            begin
//                state <= writing_to_sha;
//                writed_words_counter <= writed_words_counter + 1;
//            end
//           case(writed_words_counter_wire)
//                10'b0000010000 : state <= generating_hash;//1
//                10'b0000100000 : state <= generating_hash;//2
//                10'b0000110000 : state <= generating_hash;//3
//                10'b0001000000 : state <= final_hash_generation;//4
//                // 10'b0001010000 : state <= generating_hash;//5
//                // 10'b0001100000 : state <= generating_hash;//6
//                // 10'b0001110000 : state <= generating_hash;//7
//                // 10'b0010000000 : state <= generating_hash;//8
//                // 10'b0010010000 : state <= generating_hash;//9
//                // 10'b0010100000 : state <= generating_hash;//a
//                // 10'b0010110000 : state <= generating_hash;//b
//                // 10'b0011000000 : state <= generating_hash;//c
//                // 10'b0011010000 : state <= generating_hash;//d
//                // 10'b0011100000 : state <= generating_hash;//e
//                // 10'b0011110000 : state <= generating_hash;//f
//                // 10'b0011111111 : state <= final_hash_generation;
//                default : begin state <= writing_to_sha; end
//            endcase 
         end
         
         generating_hash: begin//przeliczania po zapisaniu 50 bloków//5
            sha3_init <= 0;
            generating_hash_counter = generating_hash_counter + 1;
            if(generating_hash_counter == 63)
            begin
                state <= hash_generated;
                generating_hash_counter <= 0; 
            end
         end
         
         hash_generated: begin///6
//            sha3_cs <= 0;
//            sha3_we <= 0;
            state <= saving_hash;//TODOdo zastanowienia
         end
         
         final_hash_generation: begin//7
            //sha3_address <= ADDR_CTRL;
            //sha3_din <= CTRL_MODE_VALUE + CTRL_INIT_VALUE;
            //sha3_cs <= 1;
            //sha3_we <= 1;
            state <= final_hash_generated ;
         end
         
         final_hash_generated: begin//8
            //sha3_cs <= 0;
            //sha3_we <= 0;
            state <= saving_hash;   
            writed_words_counter <= 0;              
         end

         saving_hash: begin//9
            case(readed_words_counter)
                4'h0 : begin sha3_address <= ADDR_DIGEST0; state <= saved_hash; end // zapisano wszystkie znaczące słowa
                4'h1 : begin sha3_address <= ADDR_DIGEST1;  state <= saved_hash; end
                4'h2 : begin sha3_address <= ADDR_DIGEST2;  state <= saved_hash; end
                4'h3 : begin sha3_address <= ADDR_DIGEST3;  state <= saved_hash; end
                4'h4 : begin sha3_address <= ADDR_DIGEST4;  state <= saved_hash; end
                4'h5 : begin sha3_address <= ADDR_DIGEST5;  state <= saved_hash; end
                4'h6 : begin sha3_address <= ADDR_DIGEST6;  state <= saved_hash; end
                4'h7 : begin sha3_address <= ADDR_DIGEST7;  state <= saved_hash; end
                4'h8 : state <= sending_data; // zapisano wszystkie znaczące słowa
                4'h9 : state <= sending_data; // zapisano wszystkie znaczące słowa
                default : sha3_address <= ADDR_DIGEST0;
            endcase
//            sha3_cs = 1;
            sha3_we = 1;
            //state <= saved_hash;
         end
         
         saved_hash: begin//10
            case(readed_words_counter)
                4'h0 : begin digest_data[31:0] <= sha3_dout; end
                4'h1 : begin digest_data[63:32] <= sha3_dout; end
                4'h2 : begin digest_data[95:64] <= sha3_dout; end
                4'h3 : begin digest_data[127:96] <= sha3_dout; end
                4'h4 : begin digest_data[159:128] <= sha3_dout; end
                4'h5 : begin digest_data[191:160] <= sha3_dout;end
                4'h6 : begin digest_data[223:192] <= sha3_dout; end
                4'h7 : begin digest_data[255:224] <= sha3_dout; end
                4'h8 : begin digest_data[287:256] <= sha3_dout; end
                4'h9 : begin digest_data[319:288] <= sha3_dout; end
                4'hA : begin digest_data[351:320] <= sha3_dout; end
                4'hB : begin digest_data[383:352] <= sha3_dout; end
                4'hC : begin digest_data[415:384] <= sha3_dout; end
                4'hD : begin digest_data[447:416] <= sha3_dout; end
                4'hE : begin digest_data[479:448] <= sha3_dout; end
                4'hF : begin digest_data[511:480] <= sha3_dout; end
                default : digest_data[31:0] <= sha3_dout;
            endcase
            sha3_we = 0;
            state <= increment_counter;
         end
         
         increment_counter : begin
            readed_words_counter = readed_words_counter + 1;
            state <= saving_hash;
         end
         
         sending_data: begin
            ready <= 1;
            case(ADDR)
                11'h000 :  DATA_OUT <= random_bits[31:0];
                11'h001 :  DATA_OUT <= random_bits[63:32];
                11'h002 :  DATA_OUT <= random_bits[95:64];
                11'h003 :  DATA_OUT <= random_bits[127:96];
                11'h004 :  DATA_OUT <= random_bits[159:128];
                11'h005 :  DATA_OUT <= random_bits[191:160];
                11'h006 :  DATA_OUT <= random_bits[223:192];
                11'h007 :  DATA_OUT <= random_bits[255:224];
                11'h008 :  DATA_OUT <= random_bits[287:256];
                11'h009 :  DATA_OUT <= random_bits[319:288];
                11'h00a :  DATA_OUT <= random_bits[351:320];
                11'h00b :  DATA_OUT <= random_bits[383:352];
                11'h00c :  DATA_OUT <= random_bits[415:384];
                11'h00d :  DATA_OUT <= random_bits[447:416];
                11'h00e :  DATA_OUT <= random_bits[479:448];
                11'h00f :  DATA_OUT <= random_bits[511:480];
                11'h010 :  DATA_OUT <= random_bits[543:512];
                11'h011 :  DATA_OUT <= random_bits[575:544];
                11'h012 :  DATA_OUT <= random_bits[607:576];
                11'h013 :  DATA_OUT <= random_bits[639:608];
                11'h014 :  DATA_OUT <= random_bits[671:640];
                11'h015 :  DATA_OUT <= random_bits[703:672];
                11'h016 :  DATA_OUT <= random_bits[735:704];
                11'h017 :  DATA_OUT <= random_bits[767:736];
                11'h018 :  DATA_OUT <= random_bits[799:768];
                11'h019 :  DATA_OUT <= random_bits[831:800];
                11'h01a :  DATA_OUT <= random_bits[863:832];
                11'h01b :  DATA_OUT <= random_bits[895:864];
                11'h01c :  DATA_OUT <= random_bits[927:896];
                11'h01d :  DATA_OUT <= random_bits[959:928];
                11'h01e :  DATA_OUT <= random_bits[991:960];
                11'h01f :  DATA_OUT <= random_bits[1023:992];
                // 11'h020 :  DATA_OUT <= random_bits[1055:1024];
                // 11'h021 :  DATA_OUT <= random_bits[1087:1056];
                // 11'h022 :  DATA_OUT <= random_bits[1119:1088];
                // 11'h023 :  DATA_OUT <= random_bits[1151:1120];
                // 11'h024 :  DATA_OUT <= random_bits[1183:1152];
                // 11'h025 :  DATA_OUT <= random_bits[1215:1184];
                // 11'h026 :  DATA_OUT <= random_bits[1247:1216];
                // 11'h027 :  DATA_OUT <= random_bits[1279:1248];
                // 11'h028 :  DATA_OUT <= random_bits[1311:1280];
                // 11'h029 :  DATA_OUT <= random_bits[1343:1312];
                // 11'h02a :  DATA_OUT <= random_bits[1375:1344];
                // 11'h02b :  DATA_OUT <= random_bits[1407:1376];
                // 11'h02c :  DATA_OUT <= random_bits[1439:1408];
                // 11'h02d :  DATA_OUT <= random_bits[1471:1440];
                // 11'h02e :  DATA_OUT <= random_bits[1503:1472];
                // 11'h02f :  DATA_OUT <= random_bits[1535:1504];
                // 11'h030 :  DATA_OUT <= random_bits[1567:1536];
                // 11'h031 :  DATA_OUT <= random_bits[1599:1568];
                // 11'h032 :  DATA_OUT <= random_bits[1631:1600];
                // 11'h033 :  DATA_OUT <= random_bits[1663:1632];
                // 11'h034 :  DATA_OUT <= random_bits[1695:1664];
                // 11'h035 :  DATA_OUT <= random_bits[1727:1696];
                // 11'h036 :  DATA_OUT <= random_bits[1759:1728];
                // 11'h037 :  DATA_OUT <= random_bits[1791:1760];
                // 11'h038 :  DATA_OUT <= random_bits[1823:1792];
                // 11'h039 :  DATA_OUT <= random_bits[1855:1824];
                // 11'h03a :  DATA_OUT <= random_bits[1887:1856];
                // 11'h03b :  DATA_OUT <= random_bits[1919:1888];
                // 11'h03c :  DATA_OUT <= random_bits[1951:1920];
                // 11'h03d :  DATA_OUT <= random_bits[1983:1952];
                // 11'h03e :  DATA_OUT <= random_bits[2015:1984];
                // 11'h03f :  DATA_OUT <= random_bits[2047:2016];
                // 11'h040 :  DATA_OUT <= random_bits[2079:2048];
                // 11'h041 :  DATA_OUT <= random_bits[2111:2080];
                // 11'h042 :  DATA_OUT <= random_bits[2143:2112];
                // 11'h043 :  DATA_OUT <= random_bits[2175:2144];
                // 11'h044 :  DATA_OUT <= random_bits[2207:2176];
                // 11'h045 :  DATA_OUT <= random_bits[2239:2208];
                // 11'h046 :  DATA_OUT <= random_bits[2271:2240];
                // 11'h047 :  DATA_OUT <= random_bits[2303:2272];
                // 11'h048 :  DATA_OUT <= random_bits[2335:2304];
                // 11'h049 :  DATA_OUT <= random_bits[2367:2336];
                // 11'h04a :  DATA_OUT <= random_bits[2399:2368];
                // 11'h04b :  DATA_OUT <= random_bits[2431:2400];
                // 11'h04c :  DATA_OUT <= random_bits[2463:2432];
                // 11'h04d :  DATA_OUT <= random_bits[2495:2464];
                // 11'h04e :  DATA_OUT <= random_bits[2527:2496];
                // 11'h04f :  DATA_OUT <= random_bits[2559:2528];
                // 11'h050 :  DATA_OUT <= random_bits[2591:2560];
                // 11'h051 :  DATA_OUT <= random_bits[2623:2592];
                // 11'h052 :  DATA_OUT <= random_bits[2655:2624];
                // 11'h053 :  DATA_OUT <= random_bits[2687:2656];
                // 11'h054 :  DATA_OUT <= random_bits[2719:2688];
                // 11'h055 :  DATA_OUT <= random_bits[2751:2720];
                // 11'h056 :  DATA_OUT <= random_bits[2783:2752];
                // 11'h057 :  DATA_OUT <= random_bits[2815:2784];
                // 11'h058 :  DATA_OUT <= random_bits[2847:2816];
                // 11'h059 :  DATA_OUT <= random_bits[2879:2848];
                // 11'h05a :  DATA_OUT <= random_bits[2911:2880];
                // 11'h05b :  DATA_OUT <= random_bits[2943:2912];
                // 11'h05c :  DATA_OUT <= random_bits[2975:2944];
                // 11'h05d :  DATA_OUT <= random_bits[3007:2976];
                // 11'h05e :  DATA_OUT <= random_bits[3039:3008];
                // 11'h05f :  DATA_OUT <= random_bits[3071:3040];
                // 11'h060 :  DATA_OUT <= random_bits[3103:3072];
                // 11'h061 :  DATA_OUT <= random_bits[3135:3104];
                // 11'h062 :  DATA_OUT <= random_bits[3167:3136];
                // 11'h063 :  DATA_OUT <= random_bits[3199:3168];
                // 11'h064 :  DATA_OUT <= random_bits[3231:3200];
                // 11'h065 :  DATA_OUT <= random_bits[3263:3232];
                // 11'h066 :  DATA_OUT <= random_bits[3295:3264];
                // 11'h067 :  DATA_OUT <= random_bits[3327:3296];
                // 11'h068 :  DATA_OUT <= random_bits[3359:3328];
                // 11'h069 :  DATA_OUT <= random_bits[3391:3360];
                // 11'h06a :  DATA_OUT <= random_bits[3423:3392];
                // 11'h06b :  DATA_OUT <= random_bits[3455:3424];
                // 11'h06c :  DATA_OUT <= random_bits[3487:3456];
                // 11'h06d :  DATA_OUT <= random_bits[3519:3488];
                // 11'h06e :  DATA_OUT <= random_bits[3551:3520];
                // 11'h06f :  DATA_OUT <= random_bits[3583:3552];
                // 11'h070 :  DATA_OUT <= random_bits[3615:3584];
                // 11'h071 :  DATA_OUT <= random_bits[3647:3616];
                // 11'h072 :  DATA_OUT <= random_bits[3679:3648];
                // 11'h073 :  DATA_OUT <= random_bits[3711:3680];
                // 11'h074 :  DATA_OUT <= random_bits[3743:3712];
                // 11'h075 :  DATA_OUT <= random_bits[3775:3744];
                // 11'h076 :  DATA_OUT <= random_bits[3807:3776];
                // 11'h077 :  DATA_OUT <= random_bits[3839:3808];
                // 11'h078 :  DATA_OUT <= random_bits[3871:3840];
                // 11'h079 :  DATA_OUT <= random_bits[3903:3872];
                // 11'h07a :  DATA_OUT <= random_bits[3935:3904];
                // 11'h07b :  DATA_OUT <= random_bits[3967:3936];
                // 11'h07c :  DATA_OUT <= random_bits[3999:3968];
                // 11'h07d :  DATA_OUT <= random_bits[4031:4000];
                // 11'h07e :  DATA_OUT <= random_bits[4063:4032];
                // 11'h07f :  DATA_OUT <= random_bits[4095:4064];
                // 11'h080 :  DATA_OUT <= random_bits[4127:4096];
                // 11'h081 :  DATA_OUT <= random_bits[4159:4128];
                // 11'h082 :  DATA_OUT <= random_bits[4191:4160];
                // 11'h083 :  DATA_OUT <= random_bits[4223:4192];
                // 11'h084 :  DATA_OUT <= random_bits[4255:4224];
                // 11'h085 :  DATA_OUT <= random_bits[4287:4256];
                // 11'h086 :  DATA_OUT <= random_bits[4319:4288];
                // 11'h087 :  DATA_OUT <= random_bits[4351:4320];
                // 11'h088 :  DATA_OUT <= random_bits[4383:4352];
                // 11'h089 :  DATA_OUT <= random_bits[4415:4384];
                // 11'h08a :  DATA_OUT <= random_bits[4447:4416];
                // 11'h08b :  DATA_OUT <= random_bits[4479:4448];
                // 11'h08c :  DATA_OUT <= random_bits[4511:4480];
                // 11'h08d :  DATA_OUT <= random_bits[4543:4512];
                // 11'h08e :  DATA_OUT <= random_bits[4575:4544];
                // 11'h08f :  DATA_OUT <= random_bits[4607:4576];
                // 11'h090 :  DATA_OUT <= random_bits[4639:4608];
                // 11'h091 :  DATA_OUT <= random_bits[4671:4640];
                // 11'h092 :  DATA_OUT <= random_bits[4703:4672];
                // 11'h093 :  DATA_OUT <= random_bits[4735:4704];
                // 11'h094 :  DATA_OUT <= random_bits[4767:4736];
                // 11'h095 :  DATA_OUT <= random_bits[4799:4768];
                // 11'h096 :  DATA_OUT <= random_bits[4831:4800];
                // 11'h097 :  DATA_OUT <= random_bits[4863:4832];
                // 11'h098 :  DATA_OUT <= random_bits[4895:4864];
                // 11'h099 :  DATA_OUT <= random_bits[4927:4896];
                // 11'h09a :  DATA_OUT <= random_bits[4959:4928];
                // 11'h09b :  DATA_OUT <= random_bits[4991:4960];
                // 11'h09c :  DATA_OUT <= random_bits[5023:4992];
                // 11'h09d :  DATA_OUT <= random_bits[5055:5024];
                // 11'h09e :  DATA_OUT <= random_bits[5087:5056];
                // 11'h09f :  DATA_OUT <= random_bits[5119:5088];
                // 11'h0a0 :  DATA_OUT <= random_bits[5151:5120];
                // 11'h0a1 :  DATA_OUT <= random_bits[5183:5152];
                // 11'h0a2 :  DATA_OUT <= random_bits[5215:5184];
                // 11'h0a3 :  DATA_OUT <= random_bits[5247:5216];
                // 11'h0a4 :  DATA_OUT <= random_bits[5279:5248];
                // 11'h0a5 :  DATA_OUT <= random_bits[5311:5280];
                // 11'h0a6 :  DATA_OUT <= random_bits[5343:5312];
                // 11'h0a7 :  DATA_OUT <= random_bits[5375:5344];
                // 11'h0a8 :  DATA_OUT <= random_bits[5407:5376];
                // 11'h0a9 :  DATA_OUT <= random_bits[5439:5408];
                // 11'h0aa :  DATA_OUT <= random_bits[5471:5440];
                // 11'h0ab :  DATA_OUT <= random_bits[5503:5472];
                // 11'h0ac :  DATA_OUT <= random_bits[5535:5504];
                // 11'h0ad :  DATA_OUT <= random_bits[5567:5536];
                // 11'h0ae :  DATA_OUT <= random_bits[5599:5568];
                // 11'h0af :  DATA_OUT <= random_bits[5631:5600];
                // 11'h0b0 :  DATA_OUT <= random_bits[5663:5632];
                // 11'h0b1 :  DATA_OUT <= random_bits[5695:5664];
                // 11'h0b2 :  DATA_OUT <= random_bits[5727:5696];
                // 11'h0b3 :  DATA_OUT <= random_bits[5759:5728];
                // 11'h0b4 :  DATA_OUT <= random_bits[5791:5760];
                // 11'h0b5 :  DATA_OUT <= random_bits[5823:5792];
                // 11'h0b6 :  DATA_OUT <= random_bits[5855:5824];
                // 11'h0b7 :  DATA_OUT <= random_bits[5887:5856];
                // 11'h0b8 :  DATA_OUT <= random_bits[5919:5888];
                // 11'h0b9 :  DATA_OUT <= random_bits[5951:5920];
                // 11'h0ba :  DATA_OUT <= random_bits[5983:5952];
                // 11'h0bb :  DATA_OUT <= random_bits[6015:5984];
                // 11'h0bc :  DATA_OUT <= random_bits[6047:6016];
                // 11'h0bd :  DATA_OUT <= random_bits[6079:6048];
                // 11'h0be :  DATA_OUT <= random_bits[6111:6080];
                // 11'h0bf :  DATA_OUT <= random_bits[6143:6112];
                // 11'h0c0 :  DATA_OUT <= random_bits[6175:6144];
                // 11'h0c1 :  DATA_OUT <= random_bits[6207:6176];
                // 11'h0c2 :  DATA_OUT <= random_bits[6239:6208];
                // 11'h0c3 :  DATA_OUT <= random_bits[6271:6240];
                // 11'h0c4 :  DATA_OUT <= random_bits[6303:6272];
                // 11'h0c5 :  DATA_OUT <= random_bits[6335:6304];
                // 11'h0c6 :  DATA_OUT <= random_bits[6367:6336];
                // 11'h0c7 :  DATA_OUT <= random_bits[6399:6368];
                // 11'h0c8 :  DATA_OUT <= random_bits[6431:6400];
                // 11'h0c9 :  DATA_OUT <= random_bits[6463:6432];
                // 11'h0ca :  DATA_OUT <= random_bits[6495:6464];
                // 11'h0cb :  DATA_OUT <= random_bits[6527:6496];
                // 11'h0cc :  DATA_OUT <= random_bits[6559:6528];
                // 11'h0cd :  DATA_OUT <= random_bits[6591:6560];
                // 11'h0ce :  DATA_OUT <= random_bits[6623:6592];
                // 11'h0cf :  DATA_OUT <= random_bits[6655:6624];
                // 11'h0d0 :  DATA_OUT <= random_bits[6687:6656];
                // 11'h0d1 :  DATA_OUT <= random_bits[6719:6688];
                // 11'h0d2 :  DATA_OUT <= random_bits[6751:6720];
                // 11'h0d3 :  DATA_OUT <= random_bits[6783:6752];
                // 11'h0d4 :  DATA_OUT <= random_bits[6815:6784];
                // 11'h0d5 :  DATA_OUT <= random_bits[6847:6816];
                // 11'h0d6 :  DATA_OUT <= random_bits[6879:6848];
                // 11'h0d7 :  DATA_OUT <= random_bits[6911:6880];
                // 11'h0d8 :  DATA_OUT <= random_bits[6943:6912];
                // 11'h0d9 :  DATA_OUT <= random_bits[6975:6944];
                // 11'h0da :  DATA_OUT <= random_bits[7007:6976];
                // 11'h0db :  DATA_OUT <= random_bits[7039:7008];
                // 11'h0dc :  DATA_OUT <= random_bits[7071:7040];
                // 11'h0dd :  DATA_OUT <= random_bits[7103:7072];
                // 11'h0de :  DATA_OUT <= random_bits[7135:7104];
                // 11'h0df :  DATA_OUT <= random_bits[7167:7136];
                // 11'h0e0 :  DATA_OUT <= random_bits[7199:7168];
                // 11'h0e1 :  DATA_OUT <= random_bits[7231:7200];
                // 11'h0e2 :  DATA_OUT <= random_bits[7263:7232];
                // 11'h0e3 :  DATA_OUT <= random_bits[7295:7264];
                // 11'h0e4 :  DATA_OUT <= random_bits[7327:7296];
                // 11'h0e5 :  DATA_OUT <= random_bits[7359:7328];
                // 11'h0e6 :  DATA_OUT <= random_bits[7391:7360];
                // 11'h0e7 :  DATA_OUT <= random_bits[7423:7392];
                // 11'h0e8 :  DATA_OUT <= random_bits[7455:7424];
                // 11'h0e9 :  DATA_OUT <= random_bits[7487:7456];
                // 11'h0ea :  DATA_OUT <= random_bits[7519:7488];
                // 11'h0eb :  DATA_OUT <= random_bits[7551:7520];
                // 11'h0ec :  DATA_OUT <= random_bits[7583:7552];
                // 11'h0ed :  DATA_OUT <= random_bits[7615:7584];
                // 11'h0ee :  DATA_OUT <= random_bits[7647:7616];
                // 11'h0ef :  DATA_OUT <= random_bits[7679:7648];
                // 11'h0f0 :  DATA_OUT <= random_bits[7711:7680];
                // 11'h0f1 :  DATA_OUT <= random_bits[7743:7712];
                // 11'h0f2 :  DATA_OUT <= random_bits[7775:7744];
                // 11'h0f3 :  DATA_OUT <= random_bits[7807:7776];
                // 11'h0f4 :  DATA_OUT <= random_bits[7839:7808];
                // 11'h0f5 :  DATA_OUT <= random_bits[7871:7840];
                // 11'h0f6 :  DATA_OUT <= random_bits[7903:7872];
                // 11'h0f7 :  DATA_OUT <= random_bits[7935:7904];
                // 11'h0f8 :  DATA_OUT <= random_bits[7967:7936];
                // 11'h0f9 :  DATA_OUT <= random_bits[7999:7968];
                // 11'h0fa :  DATA_OUT <= random_bits[8031:8000];
                // 11'h0fb :  DATA_OUT <= random_bits[8063:8032];
                // 11'h0fc :  DATA_OUT <= random_bits[8095:8064];
                // 11'h0fd :  DATA_OUT <= random_bits[8127:8096];
                // 11'h0fe :  DATA_OUT <= random_bits[8159:8128];
                // 11'h0ff :  DATA_OUT <= random_bits[8191:8160];
                // 11'h100 :  DATA_OUT <= random_bits[8223:8192];
                // 11'h101 :  DATA_OUT <= random_bits[8255:8224];
                // 11'h102 :  DATA_OUT <= random_bits[8287:8256];
                // 11'h103 :  DATA_OUT <= random_bits[8319:8288];
                // 11'h104 :  DATA_OUT <= random_bits[8351:8320];
                // 11'h105 :  DATA_OUT <= random_bits[8383:8352];
                // 11'h106 :  DATA_OUT <= random_bits[8415:8384];
                // 11'h107 :  DATA_OUT <= random_bits[8447:8416];
                // 11'h108 :  DATA_OUT <= random_bits[8479:8448];
                // 11'h109 :  DATA_OUT <= random_bits[8511:8480];
                // 11'h10a :  DATA_OUT <= random_bits[8543:8512];
                // 11'h10b :  DATA_OUT <= random_bits[8575:8544];
                // 11'h10c :  DATA_OUT <= random_bits[8607:8576];
                // 11'h10d :  DATA_OUT <= random_bits[8639:8608];
                // 11'h10e :  DATA_OUT <= random_bits[8671:8640];
                // 11'h10f :  DATA_OUT <= random_bits[8703:8672];
                // 11'h110 :  DATA_OUT <= random_bits[8735:8704];
                // 11'h111 :  DATA_OUT <= random_bits[8767:8736];
                // 11'h112 :  DATA_OUT <= random_bits[8799:8768];
                // 11'h113 :  DATA_OUT <= random_bits[8831:8800];
                // 11'h114 :  DATA_OUT <= random_bits[8863:8832];
                // 11'h115 :  DATA_OUT <= random_bits[8895:8864];
                // 11'h116 :  DATA_OUT <= random_bits[8927:8896];
                // 11'h117 :  DATA_OUT <= random_bits[8959:8928];
                // 11'h118 :  DATA_OUT <= random_bits[8991:8960];
                // 11'h119 :  DATA_OUT <= random_bits[9023:8992];
                // 11'h11a :  DATA_OUT <= random_bits[9055:9024];
                // 11'h11b :  DATA_OUT <= random_bits[9087:9056];
                // 11'h11c :  DATA_OUT <= random_bits[9119:9088];
                // 11'h11d :  DATA_OUT <= random_bits[9151:9120];
                // 11'h11e :  DATA_OUT <= random_bits[9183:9152];
                // 11'h11f :  DATA_OUT <= random_bits[9215:9184];
                // 11'h120 :  DATA_OUT <= random_bits[9247:9216];
                // 11'h121 :  DATA_OUT <= random_bits[9279:9248];
                // 11'h122 :  DATA_OUT <= random_bits[9311:9280];
                // 11'h123 :  DATA_OUT <= random_bits[9343:9312];
                // 11'h124 :  DATA_OUT <= random_bits[9375:9344];
                // 11'h125 :  DATA_OUT <= random_bits[9407:9376];
                // 11'h126 :  DATA_OUT <= random_bits[9439:9408];
                // 11'h127 :  DATA_OUT <= random_bits[9471:9440];
                // 11'h128 :  DATA_OUT <= random_bits[9503:9472];
                // 11'h129 :  DATA_OUT <= random_bits[9535:9504];
                // 11'h12a :  DATA_OUT <= random_bits[9567:9536];
                // 11'h12b :  DATA_OUT <= random_bits[9599:9568];
                // 11'h12c :  DATA_OUT <= random_bits[9631:9600];
                // 11'h12d :  DATA_OUT <= random_bits[9663:9632];
                // 11'h12e :  DATA_OUT <= random_bits[9695:9664];
                // 11'h12f :  DATA_OUT <= random_bits[9727:9696];
                // 11'h130 :  DATA_OUT <= random_bits[9759:9728];
                // 11'h131 :  DATA_OUT <= random_bits[9791:9760];
                // 11'h132 :  DATA_OUT <= random_bits[9823:9792];
                // 11'h133 :  DATA_OUT <= random_bits[9855:9824];
                // 11'h134 :  DATA_OUT <= random_bits[9887:9856];
                // 11'h135 :  DATA_OUT <= random_bits[9919:9888];
                // 11'h136 :  DATA_OUT <= random_bits[9951:9920];
                // 11'h137 :  DATA_OUT <= random_bits[9983:9952];
                // 11'h138 :  DATA_OUT <= random_bits[10015:9984];
                // 11'h139 :  DATA_OUT <= random_bits[10047:10016];
                // 11'h13a :  DATA_OUT <= random_bits[10079:10048];
                // 11'h13b :  DATA_OUT <= random_bits[10111:10080];
                // 11'h13c :  DATA_OUT <= random_bits[10143:10112];
                // 11'h13d :  DATA_OUT <= random_bits[10175:10144];
                // 11'h13e :  DATA_OUT <= random_bits[10207:10176];
                // 11'h13f :  DATA_OUT <= random_bits[10239:10208];
                // 11'h140 :  DATA_OUT <= random_bits[10271:10240];
                // 11'h141 :  DATA_OUT <= random_bits[10303:10272];
                // 11'h142 :  DATA_OUT <= random_bits[10335:10304];
                // 11'h143 :  DATA_OUT <= random_bits[10367:10336];
                // 11'h144 :  DATA_OUT <= random_bits[10399:10368];
                // 11'h145 :  DATA_OUT <= random_bits[10431:10400];
                // 11'h146 :  DATA_OUT <= random_bits[10463:10432];
                // 11'h147 :  DATA_OUT <= random_bits[10495:10464];
                // 11'h148 :  DATA_OUT <= random_bits[10527:10496];
                // 11'h149 :  DATA_OUT <= random_bits[10559:10528];
                // 11'h14a :  DATA_OUT <= random_bits[10591:10560];
                // 11'h14b :  DATA_OUT <= random_bits[10623:10592];
                // 11'h14c :  DATA_OUT <= random_bits[10655:10624];
                // 11'h14d :  DATA_OUT <= random_bits[10687:10656];
                // 11'h14e :  DATA_OUT <= random_bits[10719:10688];
                // 11'h14f :  DATA_OUT <= random_bits[10751:10720];
                // 11'h150 :  DATA_OUT <= random_bits[10783:10752];
                // 11'h151 :  DATA_OUT <= random_bits[10815:10784];
                // 11'h152 :  DATA_OUT <= random_bits[10847:10816];
                // 11'h153 :  DATA_OUT <= random_bits[10879:10848];
                // 11'h154 :  DATA_OUT <= random_bits[10911:10880];
                // 11'h155 :  DATA_OUT <= random_bits[10943:10912];
                // 11'h156 :  DATA_OUT <= random_bits[10975:10944];
                // 11'h157 :  DATA_OUT <= random_bits[11007:10976];
                // 11'h158 :  DATA_OUT <= random_bits[11039:11008];
                // 11'h159 :  DATA_OUT <= random_bits[11071:11040];
                // 11'h15a :  DATA_OUT <= random_bits[11103:11072];
                // 11'h15b :  DATA_OUT <= random_bits[11135:11104];
                // 11'h15c :  DATA_OUT <= random_bits[11167:11136];
                // 11'h15d :  DATA_OUT <= random_bits[11199:11168];
                // 11'h15e :  DATA_OUT <= random_bits[11231:11200];
                // 11'h15f :  DATA_OUT <= random_bits[11263:11232];
                // 11'h160 :  DATA_OUT <= random_bits[11295:11264];
                // 11'h161 :  DATA_OUT <= random_bits[11327:11296];
                // 11'h162 :  DATA_OUT <= random_bits[11359:11328];
                // 11'h163 :  DATA_OUT <= random_bits[11391:11360];
                // 11'h164 :  DATA_OUT <= random_bits[11423:11392];
                // 11'h165 :  DATA_OUT <= random_bits[11455:11424];
                // 11'h166 :  DATA_OUT <= random_bits[11487:11456];
                // 11'h167 :  DATA_OUT <= random_bits[11519:11488];
                // 11'h168 :  DATA_OUT <= random_bits[11551:11520];
                // 11'h169 :  DATA_OUT <= random_bits[11583:11552];
                // 11'h16a :  DATA_OUT <= random_bits[11615:11584];
                // 11'h16b :  DATA_OUT <= random_bits[11647:11616];
                // 11'h16c :  DATA_OUT <= random_bits[11679:11648];
                // 11'h16d :  DATA_OUT <= random_bits[11711:11680];
                // 11'h16e :  DATA_OUT <= random_bits[11743:11712];
                // 11'h16f :  DATA_OUT <= random_bits[11775:11744];
                // 11'h170 :  DATA_OUT <= random_bits[11807:11776];
                // 11'h171 :  DATA_OUT <= random_bits[11839:11808];
                // 11'h172 :  DATA_OUT <= random_bits[11871:11840];
                // 11'h173 :  DATA_OUT <= random_bits[11903:11872];
                // 11'h174 :  DATA_OUT <= random_bits[11935:11904];
                // 11'h175 :  DATA_OUT <= random_bits[11967:11936];
                // 11'h176 :  DATA_OUT <= random_bits[11999:11968];
                // 11'h177 :  DATA_OUT <= random_bits[12031:12000];
                // 11'h178 :  DATA_OUT <= random_bits[12063:12032];
                // 11'h179 :  DATA_OUT <= random_bits[12095:12064];
                // 11'h17a :  DATA_OUT <= random_bits[12127:12096];
                // 11'h17b :  DATA_OUT <= random_bits[12159:12128];
                // 11'h17c :  DATA_OUT <= random_bits[12191:12160];
                // 11'h17d :  DATA_OUT <= random_bits[12223:12192];
                // 11'h17e :  DATA_OUT <= random_bits[12255:12224];
                // 11'h17f :  DATA_OUT <= random_bits[12287:12256];
                // 11'h180 :  DATA_OUT <= random_bits[12319:12288];
                // 11'h181 :  DATA_OUT <= random_bits[12351:12320];
                // 11'h182 :  DATA_OUT <= random_bits[12383:12352];
                // 11'h183 :  DATA_OUT <= random_bits[12415:12384];
                // 11'h184 :  DATA_OUT <= random_bits[12447:12416];
                // 11'h185 :  DATA_OUT <= random_bits[12479:12448];
                // 11'h186 :  DATA_OUT <= random_bits[12511:12480];
                // 11'h187 :  DATA_OUT <= random_bits[12543:12512];
                // 11'h188 :  DATA_OUT <= random_bits[12575:12544];
                // 11'h189 :  DATA_OUT <= random_bits[12607:12576];
                // 11'h18a :  DATA_OUT <= random_bits[12639:12608];
                // 11'h18b :  DATA_OUT <= random_bits[12671:12640];
                // 11'h18c :  DATA_OUT <= random_bits[12703:12672];
                // 11'h18d :  DATA_OUT <= random_bits[12735:12704];
                // 11'h18e :  DATA_OUT <= random_bits[12767:12736];
                // 11'h18f :  DATA_OUT <= random_bits[12799:12768];
                // 11'h190 :  DATA_OUT <= random_bits[12831:12800];
                // 11'h191 :  DATA_OUT <= random_bits[12863:12832];
                // 11'h192 :  DATA_OUT <= random_bits[12895:12864];
                // 11'h193 :  DATA_OUT <= random_bits[12927:12896];
                // 11'h194 :  DATA_OUT <= random_bits[12959:12928];
                // 11'h195 :  DATA_OUT <= random_bits[12991:12960];
                // 11'h196 :  DATA_OUT <= random_bits[13023:12992];
                // 11'h197 :  DATA_OUT <= random_bits[13055:13024];
                // 11'h198 :  DATA_OUT <= random_bits[13087:13056];
                // 11'h199 :  DATA_OUT <= random_bits[13119:13088];
                // 11'h19a :  DATA_OUT <= random_bits[13151:13120];
                // 11'h19b :  DATA_OUT <= random_bits[13183:13152];
                // 11'h19c :  DATA_OUT <= random_bits[13215:13184];
                // 11'h19d :  DATA_OUT <= random_bits[13247:13216];
                // 11'h19e :  DATA_OUT <= random_bits[13279:13248];
                // 11'h19f :  DATA_OUT <= random_bits[13311:13280];
                // 11'h1a0 :  DATA_OUT <= random_bits[13343:13312];
                // 11'h1a1 :  DATA_OUT <= random_bits[13375:13344];
                // 11'h1a2 :  DATA_OUT <= random_bits[13407:13376];
                // 11'h1a3 :  DATA_OUT <= random_bits[13439:13408];
                // 11'h1a4 :  DATA_OUT <= random_bits[13471:13440];
                // 11'h1a5 :  DATA_OUT <= random_bits[13503:13472];
                // 11'h1a6 :  DATA_OUT <= random_bits[13535:13504];
                // 11'h1a7 :  DATA_OUT <= random_bits[13567:13536];
                // 11'h1a8 :  DATA_OUT <= random_bits[13599:13568];
                // 11'h1a9 :  DATA_OUT <= random_bits[13631:13600];
                // 11'h1aa :  DATA_OUT <= random_bits[13663:13632];
                // 11'h1ab :  DATA_OUT <= random_bits[13695:13664];
                // 11'h1ac :  DATA_OUT <= random_bits[13727:13696];
                // 11'h1ad :  DATA_OUT <= random_bits[13759:13728];
                // 11'h1ae :  DATA_OUT <= random_bits[13791:13760];
                // 11'h1af :  DATA_OUT <= random_bits[13823:13792];
                // 11'h1b0 :  DATA_OUT <= random_bits[13855:13824];
                // 11'h1b1 :  DATA_OUT <= random_bits[13887:13856];
                // 11'h1b2 :  DATA_OUT <= random_bits[13919:13888];
                // 11'h1b3 :  DATA_OUT <= random_bits[13951:13920];
                // 11'h1b4 :  DATA_OUT <= random_bits[13983:13952];
                // 11'h1b5 :  DATA_OUT <= random_bits[14015:13984];
                // 11'h1b6 :  DATA_OUT <= random_bits[14047:14016];
                // 11'h1b7 :  DATA_OUT <= random_bits[14079:14048];
                // 11'h1b8 :  DATA_OUT <= random_bits[14111:14080];
                // 11'h1b9 :  DATA_OUT <= random_bits[14143:14112];
                // 11'h1ba :  DATA_OUT <= random_bits[14175:14144];
                // 11'h1bb :  DATA_OUT <= random_bits[14207:14176];
                // 11'h1bc :  DATA_OUT <= random_bits[14239:14208];
                // 11'h1bd :  DATA_OUT <= random_bits[14271:14240];
                // 11'h1be :  DATA_OUT <= random_bits[14303:14272];
                // 11'h1bf :  DATA_OUT <= random_bits[14335:14304];
                // 11'h1c0 :  DATA_OUT <= random_bits[14367:14336];
                // 11'h1c1 :  DATA_OUT <= random_bits[14399:14368];
                // 11'h1c2 :  DATA_OUT <= random_bits[14431:14400];
                // 11'h1c3 :  DATA_OUT <= random_bits[14463:14432];
                // 11'h1c4 :  DATA_OUT <= random_bits[14495:14464];
                // 11'h1c5 :  DATA_OUT <= random_bits[14527:14496];
                // 11'h1c6 :  DATA_OUT <= random_bits[14559:14528];
                // 11'h1c7 :  DATA_OUT <= random_bits[14591:14560];
                // 11'h1c8 :  DATA_OUT <= random_bits[14623:14592];
                // 11'h1c9 :  DATA_OUT <= random_bits[14655:14624];
                // 11'h1ca :  DATA_OUT <= random_bits[14687:14656];
                // 11'h1cb :  DATA_OUT <= random_bits[14719:14688];
                // 11'h1cc :  DATA_OUT <= random_bits[14751:14720];
                // 11'h1cd :  DATA_OUT <= random_bits[14783:14752];
                // 11'h1ce :  DATA_OUT <= random_bits[14815:14784];
                // 11'h1cf :  DATA_OUT <= random_bits[14847:14816];
                // 11'h1d0 :  DATA_OUT <= random_bits[14879:14848];
                // 11'h1d1 :  DATA_OUT <= random_bits[14911:14880];
                // 11'h1d2 :  DATA_OUT <= random_bits[14943:14912];
                // 11'h1d3 :  DATA_OUT <= random_bits[14975:14944];
                // 11'h1d4 :  DATA_OUT <= random_bits[15007:14976];
                // 11'h1d5 :  DATA_OUT <= random_bits[15039:15008];
                // 11'h1d6 :  DATA_OUT <= random_bits[15071:15040];
                // 11'h1d7 :  DATA_OUT <= random_bits[15103:15072];
                // 11'h1d8 :  DATA_OUT <= random_bits[15135:15104];
                // 11'h1d9 :  DATA_OUT <= random_bits[15167:15136];
                // 11'h1da :  DATA_OUT <= random_bits[15199:15168];
                // 11'h1db :  DATA_OUT <= random_bits[15231:15200];
                // 11'h1dc :  DATA_OUT <= random_bits[15263:15232];
                // 11'h1dd :  DATA_OUT <= random_bits[15295:15264];
                // 11'h1de :  DATA_OUT <= random_bits[15327:15296];
                // 11'h1df :  DATA_OUT <= random_bits[15359:15328];
                // 11'h1e0 :  DATA_OUT <= random_bits[15391:15360];
                // 11'h1e1 :  DATA_OUT <= random_bits[15423:15392];
                // 11'h1e2 :  DATA_OUT <= random_bits[15455:15424];
                // 11'h1e3 :  DATA_OUT <= random_bits[15487:15456];
                // 11'h1e4 :  DATA_OUT <= random_bits[15519:15488];
                // 11'h1e5 :  DATA_OUT <= random_bits[15551:15520];
                // 11'h1e6 :  DATA_OUT <= random_bits[15583:15552];
                // 11'h1e7 :  DATA_OUT <= random_bits[15615:15584];
                // 11'h1e8 :  DATA_OUT <= random_bits[15647:15616];
                // 11'h1e9 :  DATA_OUT <= random_bits[15679:15648];
                // 11'h1ea :  DATA_OUT <= random_bits[15711:15680];
                // 11'h1eb :  DATA_OUT <= random_bits[15743:15712];
                // 11'h1ec :  DATA_OUT <= random_bits[15775:15744];
                // 11'h1ed :  DATA_OUT <= random_bits[15807:15776];
                // 11'h1ee :  DATA_OUT <= random_bits[15839:15808];
                // 11'h1ef :  DATA_OUT <= random_bits[15871:15840];
                // 11'h1f0 :  DATA_OUT <= random_bits[15903:15872];
                // 11'h1f1 :  DATA_OUT <= random_bits[15935:15904];
                // 11'h1f2 :  DATA_OUT <= random_bits[15967:15936];
                // 11'h1f3 :  DATA_OUT <= random_bits[15999:15968];
                // 11'h1f4 :  DATA_OUT <= random_bits[16031:16000];
                // 11'h1f5 :  DATA_OUT <= random_bits[16063:16032];
                // 11'h1f6 :  DATA_OUT <= random_bits[16095:16064];
                // 11'h1f7 :  DATA_OUT <= random_bits[16127:16096];
                // 11'h1f8 :  DATA_OUT <= random_bits[16159:16128];
                // 11'h1f9 :  DATA_OUT <= random_bits[16191:16160];
                // 11'h1fa :  DATA_OUT <= random_bits[16223:16192];
                // 11'h1fb :  DATA_OUT <= random_bits[16255:16224];
                // 11'h1fc :  DATA_OUT <= random_bits[16287:16256];
                // 11'h1fd :  DATA_OUT <= random_bits[16319:16288];
                // 11'h1fe :  DATA_OUT <= random_bits[16351:16320];
                // 11'h1ff :  DATA_OUT <= random_bits[16383:16352];
                // 11'h200 :  DATA_OUT <= random_bits[16415:16384];
                // 11'h201 :  DATA_OUT <= random_bits[16447:16416];
                // 11'h202 :  DATA_OUT <= random_bits[16479:16448];
                // 11'h203 :  DATA_OUT <= random_bits[16511:16480];
                // 11'h204 :  DATA_OUT <= random_bits[16543:16512];
                // 11'h205 :  DATA_OUT <= random_bits[16575:16544];
                // 11'h206 :  DATA_OUT <= random_bits[16607:16576];
                // 11'h207 :  DATA_OUT <= random_bits[16639:16608];
                // 11'h208 :  DATA_OUT <= random_bits[16671:16640];
                // 11'h209 :  DATA_OUT <= random_bits[16703:16672];
                // 11'h20a :  DATA_OUT <= random_bits[16735:16704];
                // 11'h20b :  DATA_OUT <= random_bits[16767:16736];
                // 11'h20c :  DATA_OUT <= random_bits[16799:16768];
                // 11'h20d :  DATA_OUT <= random_bits[16831:16800];
                // 11'h20e :  DATA_OUT <= random_bits[16863:16832];
                // 11'h20f :  DATA_OUT <= random_bits[16895:16864];
                // 11'h210 :  DATA_OUT <= random_bits[16927:16896];
                // 11'h211 :  DATA_OUT <= random_bits[16959:16928];
                // 11'h212 :  DATA_OUT <= random_bits[16991:16960];
                // 11'h213 :  DATA_OUT <= random_bits[17023:16992];
                // 11'h214 :  DATA_OUT <= random_bits[17055:17024];
                // 11'h215 :  DATA_OUT <= random_bits[17087:17056];
                // 11'h216 :  DATA_OUT <= random_bits[17119:17088];
                // 11'h217 :  DATA_OUT <= random_bits[17151:17120];
                // 11'h218 :  DATA_OUT <= random_bits[17183:17152];
                // 11'h219 :  DATA_OUT <= random_bits[17215:17184];
                // 11'h21a :  DATA_OUT <= random_bits[17247:17216];
                // 11'h21b :  DATA_OUT <= random_bits[17279:17248];
                // 11'h21c :  DATA_OUT <= random_bits[17311:17280];
                // 11'h21d :  DATA_OUT <= random_bits[17343:17312];
                // 11'h21e :  DATA_OUT <= random_bits[17375:17344];
                // 11'h21f :  DATA_OUT <= random_bits[17407:17376];
                // 11'h220 :  DATA_OUT <= random_bits[17439:17408];
                // 11'h221 :  DATA_OUT <= random_bits[17471:17440];
                // 11'h222 :  DATA_OUT <= random_bits[17503:17472];
                // 11'h223 :  DATA_OUT <= random_bits[17535:17504];
                // 11'h224 :  DATA_OUT <= random_bits[17567:17536];
                // 11'h225 :  DATA_OUT <= random_bits[17599:17568];
                // 11'h226 :  DATA_OUT <= random_bits[17631:17600];
                // 11'h227 :  DATA_OUT <= random_bits[17663:17632];
                // 11'h228 :  DATA_OUT <= random_bits[17695:17664];
                // 11'h229 :  DATA_OUT <= random_bits[17727:17696];
                // 11'h22a :  DATA_OUT <= random_bits[17759:17728];
                // 11'h22b :  DATA_OUT <= random_bits[17791:17760];
                // 11'h22c :  DATA_OUT <= random_bits[17823:17792];
                // 11'h22d :  DATA_OUT <= random_bits[17855:17824];
                // 11'h22e :  DATA_OUT <= random_bits[17887:17856];
                // 11'h22f :  DATA_OUT <= random_bits[17919:17888];
                // 11'h230 :  DATA_OUT <= random_bits[17951:17920];
                // 11'h231 :  DATA_OUT <= random_bits[17983:17952];
                // 11'h232 :  DATA_OUT <= random_bits[18015:17984];
                // 11'h233 :  DATA_OUT <= random_bits[18047:18016];
                // 11'h234 :  DATA_OUT <= random_bits[18079:18048];
                // 11'h235 :  DATA_OUT <= random_bits[18111:18080];
                // 11'h236 :  DATA_OUT <= random_bits[18143:18112];
                // 11'h237 :  DATA_OUT <= random_bits[18175:18144];
                // 11'h238 :  DATA_OUT <= random_bits[18207:18176];
                // 11'h239 :  DATA_OUT <= random_bits[18239:18208];
                // 11'h23a :  DATA_OUT <= random_bits[18271:18240];
                // 11'h23b :  DATA_OUT <= random_bits[18303:18272];
                // 11'h23c :  DATA_OUT <= random_bits[18335:18304];
                // 11'h23d :  DATA_OUT <= random_bits[18367:18336];
                // 11'h23e :  DATA_OUT <= random_bits[18399:18368];
                // 11'h23f :  DATA_OUT <= random_bits[18431:18400];
                // 11'h240 :  DATA_OUT <= random_bits[18463:18432];
                // 11'h241 :  DATA_OUT <= random_bits[18495:18464];
                // 11'h242 :  DATA_OUT <= random_bits[18527:18496];
                // 11'h243 :  DATA_OUT <= random_bits[18559:18528];
                // 11'h244 :  DATA_OUT <= random_bits[18591:18560];
                // 11'h245 :  DATA_OUT <= random_bits[18623:18592];
                // 11'h246 :  DATA_OUT <= random_bits[18655:18624];
                // 11'h247 :  DATA_OUT <= random_bits[18687:18656];
                // 11'h248 :  DATA_OUT <= random_bits[18719:18688];
                // 11'h249 :  DATA_OUT <= random_bits[18751:18720];
                // 11'h24a :  DATA_OUT <= random_bits[18783:18752];
                // 11'h24b :  DATA_OUT <= random_bits[18815:18784];
                // 11'h24c :  DATA_OUT <= random_bits[18847:18816];
                // 11'h24d :  DATA_OUT <= random_bits[18879:18848];
                // 11'h24e :  DATA_OUT <= random_bits[18911:18880];
                // 11'h24f :  DATA_OUT <= random_bits[18943:18912];
                // 11'h250 :  DATA_OUT <= random_bits[18975:18944];
                // 11'h251 :  DATA_OUT <= random_bits[19007:18976];
                // 11'h252 :  DATA_OUT <= random_bits[19039:19008];
                // 11'h253 :  DATA_OUT <= random_bits[19071:19040];
                // 11'h254 :  DATA_OUT <= random_bits[19103:19072];
                // 11'h255 :  DATA_OUT <= random_bits[19135:19104];
                // 11'h256 :  DATA_OUT <= random_bits[19167:19136];
                // 11'h257 :  DATA_OUT <= random_bits[19199:19168];
                // 11'h258 :  DATA_OUT <= random_bits[19231:19200];
                // 11'h259 :  DATA_OUT <= random_bits[19263:19232];
                // 11'h25a :  DATA_OUT <= random_bits[19295:19264];
                // 11'h25b :  DATA_OUT <= random_bits[19327:19296];
                // 11'h25c :  DATA_OUT <= random_bits[19359:19328];
                // 11'h25d :  DATA_OUT <= random_bits[19391:19360];
                // 11'h25e :  DATA_OUT <= random_bits[19423:19392];
                // 11'h25f :  DATA_OUT <= random_bits[19455:19424];
                // 11'h260 :  DATA_OUT <= random_bits[19487:19456];
                // 11'h261 :  DATA_OUT <= random_bits[19519:19488];
                // 11'h262 :  DATA_OUT <= random_bits[19551:19520];
                // 11'h263 :  DATA_OUT <= random_bits[19583:19552];
                // 11'h264 :  DATA_OUT <= random_bits[19615:19584];
                // 11'h265 :  DATA_OUT <= random_bits[19647:19616];
                // 11'h266 :  DATA_OUT <= random_bits[19679:19648];
                // 11'h267 :  DATA_OUT <= random_bits[19711:19680];
                // 11'h268 :  DATA_OUT <= random_bits[19743:19712];
                // 11'h269 :  DATA_OUT <= random_bits[19775:19744];
                // 11'h26a :  DATA_OUT <= random_bits[19807:19776];
                // 11'h26b :  DATA_OUT <= random_bits[19839:19808];
                // 11'h26c :  DATA_OUT <= random_bits[19871:19840];
                // 11'h26d :  DATA_OUT <= random_bits[19903:19872];
                // 11'h26e :  DATA_OUT <= random_bits[19935:19904];
                // 11'h26f :  DATA_OUT <= random_bits[19967:19936];
                // 11'h270 :  DATA_OUT <= random_bits[19999:19968];
                // 11'h271 :  DATA_OUT <= random_bits[20031:20000];
                // 11'h272 :  DATA_OUT <= random_bits[20063:20032];
                // 11'h273 :  DATA_OUT <= random_bits[20095:20064];
                // 11'h274 :  DATA_OUT <= random_bits[20127:20096];
                // 11'h275 :  DATA_OUT <= random_bits[20159:20128];
                // 11'h276 :  DATA_OUT <= random_bits[20191:20160];
                // 11'h277 :  DATA_OUT <= random_bits[20223:20192];
                // 11'h278 :  DATA_OUT <= random_bits[20255:20224];
                // 11'h279 :  DATA_OUT <= random_bits[20287:20256];
                // 11'h27a :  DATA_OUT <= random_bits[20319:20288];
                // 11'h27b :  DATA_OUT <= random_bits[20351:20320];
                // 11'h27c :  DATA_OUT <= random_bits[20383:20352];
                // 11'h27d :  DATA_OUT <= random_bits[20415:20384];
                // 11'h27e :  DATA_OUT <= random_bits[20447:20416];
                // 11'h27f :  DATA_OUT <= random_bits[20479:20448];
                // 11'h280 :  DATA_OUT <= random_bits[20511:20480];
                // 11'h281 :  DATA_OUT <= random_bits[20543:20512];
                // 11'h282 :  DATA_OUT <= random_bits[20575:20544];
                // 11'h283 :  DATA_OUT <= random_bits[20607:20576];
                // 11'h284 :  DATA_OUT <= random_bits[20639:20608];
                // 11'h285 :  DATA_OUT <= random_bits[20671:20640];
                // 11'h286 :  DATA_OUT <= random_bits[20703:20672];
                // 11'h287 :  DATA_OUT <= random_bits[20735:20704];
                // 11'h288 :  DATA_OUT <= random_bits[20767:20736];
                // 11'h289 :  DATA_OUT <= random_bits[20799:20768];
                // 11'h28a :  DATA_OUT <= random_bits[20831:20800];
                // 11'h28b :  DATA_OUT <= random_bits[20863:20832];
                // 11'h28c :  DATA_OUT <= random_bits[20895:20864];
                // 11'h28d :  DATA_OUT <= random_bits[20927:20896];
                // 11'h28e :  DATA_OUT <= random_bits[20959:20928];
                // 11'h28f :  DATA_OUT <= random_bits[20991:20960];
                // 11'h290 :  DATA_OUT <= random_bits[21023:20992];
                // 11'h291 :  DATA_OUT <= random_bits[21055:21024];
                // 11'h292 :  DATA_OUT <= random_bits[21087:21056];
                // 11'h293 :  DATA_OUT <= random_bits[21119:21088];
                // 11'h294 :  DATA_OUT <= random_bits[21151:21120];
                // 11'h295 :  DATA_OUT <= random_bits[21183:21152];
                // 11'h296 :  DATA_OUT <= random_bits[21215:21184];
                // 11'h297 :  DATA_OUT <= random_bits[21247:21216];
                // 11'h298 :  DATA_OUT <= random_bits[21279:21248];
                // 11'h299 :  DATA_OUT <= random_bits[21311:21280];
                // 11'h29a :  DATA_OUT <= random_bits[21343:21312];
                // 11'h29b :  DATA_OUT <= random_bits[21375:21344];
                // 11'h29c :  DATA_OUT <= random_bits[21407:21376];
                // 11'h29d :  DATA_OUT <= random_bits[21439:21408];
                // 11'h29e :  DATA_OUT <= random_bits[21471:21440];
                // 11'h29f :  DATA_OUT <= random_bits[21503:21472];
                // 11'h2a0 :  DATA_OUT <= random_bits[21535:21504];
                // 11'h2a1 :  DATA_OUT <= random_bits[21567:21536];
                // 11'h2a2 :  DATA_OUT <= random_bits[21599:21568];
                // 11'h2a3 :  DATA_OUT <= random_bits[21631:21600];
                // 11'h2a4 :  DATA_OUT <= random_bits[21663:21632];
                // 11'h2a5 :  DATA_OUT <= random_bits[21695:21664];
                // 11'h2a6 :  DATA_OUT <= random_bits[21727:21696];
                // 11'h2a7 :  DATA_OUT <= random_bits[21759:21728];
                // 11'h2a8 :  DATA_OUT <= random_bits[21791:21760];
                // 11'h2a9 :  DATA_OUT <= random_bits[21823:21792];
                // 11'h2aa :  DATA_OUT <= random_bits[21855:21824];
                // 11'h2ab :  DATA_OUT <= random_bits[21887:21856];
                // 11'h2ac :  DATA_OUT <= random_bits[21919:21888];
                // 11'h2ad :  DATA_OUT <= random_bits[21951:21920];
                // 11'h2ae :  DATA_OUT <= random_bits[21983:21952];
                // 11'h2af :  DATA_OUT <= random_bits[22015:21984];
                // 11'h2b0 :  DATA_OUT <= random_bits[22047:22016];
                // 11'h2b1 :  DATA_OUT <= random_bits[22079:22048];
                // 11'h2b2 :  DATA_OUT <= random_bits[22111:22080];
                // 11'h2b3 :  DATA_OUT <= random_bits[22143:22112];
                // 11'h2b4 :  DATA_OUT <= random_bits[22175:22144];
                // 11'h2b5 :  DATA_OUT <= random_bits[22207:22176];
                // 11'h2b6 :  DATA_OUT <= random_bits[22239:22208];
                // 11'h2b7 :  DATA_OUT <= random_bits[22271:22240];
                // 11'h2b8 :  DATA_OUT <= random_bits[22303:22272];
                // 11'h2b9 :  DATA_OUT <= random_bits[22335:22304];
                // 11'h2ba :  DATA_OUT <= random_bits[22367:22336];
                // 11'h2bb :  DATA_OUT <= random_bits[22399:22368];
                // 11'h2bc :  DATA_OUT <= random_bits[22431:22400];
                // 11'h2bd :  DATA_OUT <= random_bits[22463:22432];
                // 11'h2be :  DATA_OUT <= random_bits[22495:22464];
                // 11'h2bf :  DATA_OUT <= random_bits[22527:22496];
                // 11'h2c0 :  DATA_OUT <= random_bits[22559:22528];
                // 11'h2c1 :  DATA_OUT <= random_bits[22591:22560];
                // 11'h2c2 :  DATA_OUT <= random_bits[22623:22592];
                // 11'h2c3 :  DATA_OUT <= random_bits[22655:22624];
                // 11'h2c4 :  DATA_OUT <= random_bits[22687:22656];
                // 11'h2c5 :  DATA_OUT <= random_bits[22719:22688];
                // 11'h2c6 :  DATA_OUT <= random_bits[22751:22720];
                // 11'h2c7 :  DATA_OUT <= random_bits[22783:22752];
                // 11'h2c8 :  DATA_OUT <= random_bits[22815:22784];
                // 11'h2c9 :  DATA_OUT <= random_bits[22847:22816];
                // 11'h2ca :  DATA_OUT <= random_bits[22879:22848];
                // 11'h2cb :  DATA_OUT <= random_bits[22911:22880];
                // 11'h2cc :  DATA_OUT <= random_bits[22943:22912];
                // 11'h2cd :  DATA_OUT <= random_bits[22975:22944];
                // 11'h2ce :  DATA_OUT <= random_bits[23007:22976];
                // 11'h2cf :  DATA_OUT <= random_bits[23039:23008];
                // 11'h2d0 :  DATA_OUT <= random_bits[23071:23040];
                // 11'h2d1 :  DATA_OUT <= random_bits[23103:23072];
                // 11'h2d2 :  DATA_OUT <= random_bits[23135:23104];
                // 11'h2d3 :  DATA_OUT <= random_bits[23167:23136];
                // 11'h2d4 :  DATA_OUT <= random_bits[23199:23168];
                // 11'h2d5 :  DATA_OUT <= random_bits[23231:23200];
                // 11'h2d6 :  DATA_OUT <= random_bits[23263:23232];
                // 11'h2d7 :  DATA_OUT <= random_bits[23295:23264];
                // 11'h2d8 :  DATA_OUT <= random_bits[23327:23296];
                // 11'h2d9 :  DATA_OUT <= random_bits[23359:23328];
                // 11'h2da :  DATA_OUT <= random_bits[23391:23360];
                // 11'h2db :  DATA_OUT <= random_bits[23423:23392];
                // 11'h2dc :  DATA_OUT <= random_bits[23455:23424];
                // 11'h2dd :  DATA_OUT <= random_bits[23487:23456];
                // 11'h2de :  DATA_OUT <= random_bits[23519:23488];
                // 11'h2df :  DATA_OUT <= random_bits[23551:23520];
                // 11'h2e0 :  DATA_OUT <= random_bits[23583:23552];
                // 11'h2e1 :  DATA_OUT <= random_bits[23615:23584];
                // 11'h2e2 :  DATA_OUT <= random_bits[23647:23616];
                // 11'h2e3 :  DATA_OUT <= random_bits[23679:23648];
                // 11'h2e4 :  DATA_OUT <= random_bits[23711:23680];
                // 11'h2e5 :  DATA_OUT <= random_bits[23743:23712];
                // 11'h2e6 :  DATA_OUT <= random_bits[23775:23744];
                // 11'h2e7 :  DATA_OUT <= random_bits[23807:23776];
                // 11'h2e8 :  DATA_OUT <= random_bits[23839:23808];
                // 11'h2e9 :  DATA_OUT <= random_bits[23871:23840];
                // 11'h2ea :  DATA_OUT <= random_bits[23903:23872];
                // 11'h2eb :  DATA_OUT <= random_bits[23935:23904];
                // 11'h2ec :  DATA_OUT <= random_bits[23967:23936];
                // 11'h2ed :  DATA_OUT <= random_bits[23999:23968];
                // 11'h2ee :  DATA_OUT <= random_bits[24031:24000];
                // 11'h2ef :  DATA_OUT <= random_bits[24063:24032];
                // 11'h2f0 :  DATA_OUT <= random_bits[24095:24064];
                // 11'h2f1 :  DATA_OUT <= random_bits[24127:24096];
                // 11'h2f2 :  DATA_OUT <= random_bits[24159:24128];
                // 11'h2f3 :  DATA_OUT <= random_bits[24191:24160];
                // 11'h2f4 :  DATA_OUT <= random_bits[24223:24192];
                // 11'h2f5 :  DATA_OUT <= random_bits[24255:24224];
                // 11'h2f6 :  DATA_OUT <= random_bits[24287:24256];
                // 11'h2f7 :  DATA_OUT <= random_bits[24319:24288];
                // 11'h2f8 :  DATA_OUT <= random_bits[24351:24320];
                // 11'h2f9 :  DATA_OUT <= random_bits[24383:24352];
                // 11'h2fa :  DATA_OUT <= random_bits[24415:24384];
                // 11'h2fb :  DATA_OUT <= random_bits[24447:24416];
                // 11'h2fc :  DATA_OUT <= random_bits[24479:24448];
                // 11'h2fd :  DATA_OUT <= random_bits[24511:24480];
                // 11'h2fe :  DATA_OUT <= random_bits[24543:24512];
                // 11'h2ff :  DATA_OUT <= random_bits[24575:24544];
                // 11'h300 :  DATA_OUT <= random_bits[24607:24576];
                // 11'h301 :  DATA_OUT <= random_bits[24639:24608];
                // 11'h302 :  DATA_OUT <= random_bits[24671:24640];
                // 11'h303 :  DATA_OUT <= random_bits[24703:24672];
                // 11'h304 :  DATA_OUT <= random_bits[24735:24704];
                // 11'h305 :  DATA_OUT <= random_bits[24767:24736];
                // 11'h306 :  DATA_OUT <= random_bits[24799:24768];
                // 11'h307 :  DATA_OUT <= random_bits[24831:24800];
                // 11'h308 :  DATA_OUT <= random_bits[24863:24832];
                // 11'h309 :  DATA_OUT <= random_bits[24895:24864];
                // 11'h30a :  DATA_OUT <= random_bits[24927:24896];
                // 11'h30b :  DATA_OUT <= random_bits[24959:24928];
                // 11'h30c :  DATA_OUT <= random_bits[24991:24960];
                // 11'h30d :  DATA_OUT <= random_bits[25023:24992];
                // 11'h30e :  DATA_OUT <= random_bits[25055:25024];
                // 11'h30f :  DATA_OUT <= random_bits[25087:25056];
                // 11'h310 :  DATA_OUT <= random_bits[25119:25088];
                // 11'h311 :  DATA_OUT <= random_bits[25151:25120];
                // 11'h312 :  DATA_OUT <= random_bits[25183:25152];
                // 11'h313 :  DATA_OUT <= random_bits[25215:25184];
                // 11'h314 :  DATA_OUT <= random_bits[25247:25216];
                // 11'h315 :  DATA_OUT <= random_bits[25279:25248];
                // 11'h316 :  DATA_OUT <= random_bits[25311:25280];
                // 11'h317 :  DATA_OUT <= random_bits[25343:25312];
                // 11'h318 :  DATA_OUT <= random_bits[25375:25344];
                // 11'h319 :  DATA_OUT <= random_bits[25407:25376];
                // 11'h31a :  DATA_OUT <= random_bits[25439:25408];
                // 11'h31b :  DATA_OUT <= random_bits[25471:25440];
                // 11'h31c :  DATA_OUT <= random_bits[25503:25472];
                // 11'h31d :  DATA_OUT <= random_bits[25535:25504];
                // 11'h31e :  DATA_OUT <= random_bits[25567:25536];
                // 11'h31f :  DATA_OUT <= random_bits[25599:25568];
                // 11'h320 :  DATA_OUT <= random_bits[25631:25600];
                // 11'h321 :  DATA_OUT <= random_bits[25663:25632];
                // 11'h322 :  DATA_OUT <= random_bits[25695:25664];
                // 11'h323 :  DATA_OUT <= random_bits[25727:25696];
                // 11'h324 :  DATA_OUT <= random_bits[25759:25728];
                // 11'h325 :  DATA_OUT <= random_bits[25791:25760];
                // 11'h326 :  DATA_OUT <= random_bits[25823:25792];
                // 11'h327 :  DATA_OUT <= random_bits[25855:25824];
                // 11'h328 :  DATA_OUT <= random_bits[25887:25856];
                // 11'h329 :  DATA_OUT <= random_bits[25919:25888];
                // 11'h32a :  DATA_OUT <= random_bits[25951:25920];
                // 11'h32b :  DATA_OUT <= random_bits[25983:25952];
                // 11'h32c :  DATA_OUT <= random_bits[26015:25984];
                // 11'h32d :  DATA_OUT <= random_bits[26047:26016];
                // 11'h32e :  DATA_OUT <= random_bits[26079:26048];
                // 11'h32f :  DATA_OUT <= random_bits[26111:26080];
                // 11'h330 :  DATA_OUT <= random_bits[26143:26112];
                // 11'h331 :  DATA_OUT <= random_bits[26175:26144];
                // 11'h332 :  DATA_OUT <= random_bits[26207:26176];
                // 11'h333 :  DATA_OUT <= random_bits[26239:26208];
                // 11'h334 :  DATA_OUT <= random_bits[26271:26240];
                // 11'h335 :  DATA_OUT <= random_bits[26303:26272];
                // 11'h336 :  DATA_OUT <= random_bits[26335:26304];
                // 11'h337 :  DATA_OUT <= random_bits[26367:26336];
                // 11'h338 :  DATA_OUT <= random_bits[26399:26368];
                // 11'h339 :  DATA_OUT <= random_bits[26431:26400];
                // 11'h33a :  DATA_OUT <= random_bits[26463:26432];
                // 11'h33b :  DATA_OUT <= random_bits[26495:26464];
                // 11'h33c :  DATA_OUT <= random_bits[26527:26496];
                // 11'h33d :  DATA_OUT <= random_bits[26559:26528];
                // 11'h33e :  DATA_OUT <= random_bits[26591:26560];
                // 11'h33f :  DATA_OUT <= random_bits[26623:26592];
                // 11'h340 :  DATA_OUT <= random_bits[26655:26624];
                // 11'h341 :  DATA_OUT <= random_bits[26687:26656];
                // 11'h342 :  DATA_OUT <= random_bits[26719:26688];
                // 11'h343 :  DATA_OUT <= random_bits[26751:26720];
                // 11'h344 :  DATA_OUT <= random_bits[26783:26752];
                // 11'h345 :  DATA_OUT <= random_bits[26815:26784];
                // 11'h346 :  DATA_OUT <= random_bits[26847:26816];
                // 11'h347 :  DATA_OUT <= random_bits[26879:26848];
                // 11'h348 :  DATA_OUT <= random_bits[26911:26880];
                // 11'h349 :  DATA_OUT <= random_bits[26943:26912];
                // 11'h34a :  DATA_OUT <= random_bits[26975:26944];
                // 11'h34b :  DATA_OUT <= random_bits[27007:26976];
                // 11'h34c :  DATA_OUT <= random_bits[27039:27008];
                // 11'h34d :  DATA_OUT <= random_bits[27071:27040];
                // 11'h34e :  DATA_OUT <= random_bits[27103:27072];
                // 11'h34f :  DATA_OUT <= random_bits[27135:27104];
                // 11'h350 :  DATA_OUT <= random_bits[27167:27136];
                // 11'h351 :  DATA_OUT <= random_bits[27199:27168];
                // 11'h352 :  DATA_OUT <= random_bits[27231:27200];
                // 11'h353 :  DATA_OUT <= random_bits[27263:27232];
                // 11'h354 :  DATA_OUT <= random_bits[27295:27264];
                // 11'h355 :  DATA_OUT <= random_bits[27327:27296];
                // 11'h356 :  DATA_OUT <= random_bits[27359:27328];
                // 11'h357 :  DATA_OUT <= random_bits[27391:27360];
                // 11'h358 :  DATA_OUT <= random_bits[27423:27392];
                // 11'h359 :  DATA_OUT <= random_bits[27455:27424];
                // 11'h35a :  DATA_OUT <= random_bits[27487:27456];
                // 11'h35b :  DATA_OUT <= random_bits[27519:27488];
                // 11'h35c :  DATA_OUT <= random_bits[27551:27520];
                // 11'h35d :  DATA_OUT <= random_bits[27583:27552];
                // 11'h35e :  DATA_OUT <= random_bits[27615:27584];
                // 11'h35f :  DATA_OUT <= random_bits[27647:27616];
                // 11'h360 :  DATA_OUT <= random_bits[27679:27648];
                // 11'h361 :  DATA_OUT <= random_bits[27711:27680];
                // 11'h362 :  DATA_OUT <= random_bits[27743:27712];
                // 11'h363 :  DATA_OUT <= random_bits[27775:27744];
                // 11'h364 :  DATA_OUT <= random_bits[27807:27776];
                // 11'h365 :  DATA_OUT <= random_bits[27839:27808];
                // 11'h366 :  DATA_OUT <= random_bits[27871:27840];
                // 11'h367 :  DATA_OUT <= random_bits[27903:27872];
                // 11'h368 :  DATA_OUT <= random_bits[27935:27904];
                // 11'h369 :  DATA_OUT <= random_bits[27967:27936];
                // 11'h36a :  DATA_OUT <= random_bits[27999:27968];
                // 11'h36b :  DATA_OUT <= random_bits[28031:28000];
                // 11'h36c :  DATA_OUT <= random_bits[28063:28032];
                // 11'h36d :  DATA_OUT <= random_bits[28095:28064];
                // 11'h36e :  DATA_OUT <= random_bits[28127:28096];
                // 11'h36f :  DATA_OUT <= random_bits[28159:28128];
                // 11'h370 :  DATA_OUT <= random_bits[28191:28160];
                // 11'h371 :  DATA_OUT <= random_bits[28223:28192];
                // 11'h372 :  DATA_OUT <= random_bits[28255:28224];
                // 11'h373 :  DATA_OUT <= random_bits[28287:28256];
                // 11'h374 :  DATA_OUT <= random_bits[28319:28288];
                // 11'h375 :  DATA_OUT <= random_bits[28351:28320];
                // 11'h376 :  DATA_OUT <= random_bits[28383:28352];
                // 11'h377 :  DATA_OUT <= random_bits[28415:28384];
                // 11'h378 :  DATA_OUT <= random_bits[28447:28416];
                // 11'h379 :  DATA_OUT <= random_bits[28479:28448];
                // 11'h37a :  DATA_OUT <= random_bits[28511:28480];
                // 11'h37b :  DATA_OUT <= random_bits[28543:28512];
                // 11'h37c :  DATA_OUT <= random_bits[28575:28544];
                // 11'h37d :  DATA_OUT <= random_bits[28607:28576];
                // 11'h37e :  DATA_OUT <= random_bits[28639:28608];
                // 11'h37f :  DATA_OUT <= random_bits[28671:28640];
                // 11'h380 :  DATA_OUT <= random_bits[28703:28672];
                // 11'h381 :  DATA_OUT <= random_bits[28735:28704];
                // 11'h382 :  DATA_OUT <= random_bits[28767:28736];
                // 11'h383 :  DATA_OUT <= random_bits[28799:28768];
                // 11'h384 :  DATA_OUT <= random_bits[28831:28800];
                // 11'h385 :  DATA_OUT <= random_bits[28863:28832];
                // 11'h386 :  DATA_OUT <= random_bits[28895:28864];
                // 11'h387 :  DATA_OUT <= random_bits[28927:28896];
                // 11'h388 :  DATA_OUT <= random_bits[28959:28928];
                // 11'h389 :  DATA_OUT <= random_bits[28991:28960];
                // 11'h38a :  DATA_OUT <= random_bits[29023:28992];
                // 11'h38b :  DATA_OUT <= random_bits[29055:29024];
                // 11'h38c :  DATA_OUT <= random_bits[29087:29056];
                // 11'h38d :  DATA_OUT <= random_bits[29119:29088];
                // 11'h38e :  DATA_OUT <= random_bits[29151:29120];
                // 11'h38f :  DATA_OUT <= random_bits[29183:29152];
                // 11'h390 :  DATA_OUT <= random_bits[29215:29184];
                // 11'h391 :  DATA_OUT <= random_bits[29247:29216];
                // 11'h392 :  DATA_OUT <= random_bits[29279:29248];
                // 11'h393 :  DATA_OUT <= random_bits[29311:29280];
                // 11'h394 :  DATA_OUT <= random_bits[29343:29312];
                // 11'h395 :  DATA_OUT <= random_bits[29375:29344];
                // 11'h396 :  DATA_OUT <= random_bits[29407:29376];
                // 11'h397 :  DATA_OUT <= random_bits[29439:29408];
                // 11'h398 :  DATA_OUT <= random_bits[29471:29440];
                // 11'h399 :  DATA_OUT <= random_bits[29503:29472];
                // 11'h39a :  DATA_OUT <= random_bits[29535:29504];
                // 11'h39b :  DATA_OUT <= random_bits[29567:29536];
                // 11'h39c :  DATA_OUT <= random_bits[29599:29568];
                // 11'h39d :  DATA_OUT <= random_bits[29631:29600];
                // 11'h39e :  DATA_OUT <= random_bits[29663:29632];
                // 11'h39f :  DATA_OUT <= random_bits[29695:29664];
                // 11'h3a0 :  DATA_OUT <= random_bits[29727:29696];
                // 11'h3a1 :  DATA_OUT <= random_bits[29759:29728];
                // 11'h3a2 :  DATA_OUT <= random_bits[29791:29760];
                // 11'h3a3 :  DATA_OUT <= random_bits[29823:29792];
                // 11'h3a4 :  DATA_OUT <= random_bits[29855:29824];
                // 11'h3a5 :  DATA_OUT <= random_bits[29887:29856];
                // 11'h3a6 :  DATA_OUT <= random_bits[29919:29888];
                // 11'h3a7 :  DATA_OUT <= random_bits[29951:29920];
                // 11'h3a8 :  DATA_OUT <= random_bits[29983:29952];
                // 11'h3a9 :  DATA_OUT <= random_bits[30015:29984];
                // 11'h3aa :  DATA_OUT <= random_bits[30047:30016];
                // 11'h3ab :  DATA_OUT <= random_bits[30079:30048];
                // 11'h3ac :  DATA_OUT <= random_bits[30111:30080];
                // 11'h3ad :  DATA_OUT <= random_bits[30143:30112];
                // 11'h3ae :  DATA_OUT <= random_bits[30175:30144];
                // 11'h3af :  DATA_OUT <= random_bits[30207:30176];
                // 11'h3b0 :  DATA_OUT <= random_bits[30239:30208];
                // 11'h3b1 :  DATA_OUT <= random_bits[30271:30240];
                // 11'h3b2 :  DATA_OUT <= random_bits[30303:30272];
                // 11'h3b3 :  DATA_OUT <= random_bits[30335:30304];
                // 11'h3b4 :  DATA_OUT <= random_bits[30367:30336];
                // 11'h3b5 :  DATA_OUT <= random_bits[30399:30368];
                // 11'h3b6 :  DATA_OUT <= random_bits[30431:30400];
                // 11'h3b7 :  DATA_OUT <= random_bits[30463:30432];
                // 11'h3b8 :  DATA_OUT <= random_bits[30495:30464];
                // 11'h3b9 :  DATA_OUT <= random_bits[30527:30496];
                // 11'h3ba :  DATA_OUT <= random_bits[30559:30528];
                // 11'h3bb :  DATA_OUT <= random_bits[30591:30560];
                // 11'h3bc :  DATA_OUT <= random_bits[30623:30592];
                // 11'h3bd :  DATA_OUT <= random_bits[30655:30624];
                // 11'h3be :  DATA_OUT <= random_bits[30687:30656];
                // 11'h3bf :  DATA_OUT <= random_bits[30719:30688];
                // 11'h3c0 :  DATA_OUT <= random_bits[30751:30720];
                // 11'h3c1 :  DATA_OUT <= random_bits[30783:30752];
                // 11'h3c2 :  DATA_OUT <= random_bits[30815:30784];
                // 11'h3c3 :  DATA_OUT <= random_bits[30847:30816];
                // 11'h3c4 :  DATA_OUT <= random_bits[30879:30848];
                // 11'h3c5 :  DATA_OUT <= random_bits[30911:30880];
                // 11'h3c6 :  DATA_OUT <= random_bits[30943:30912];
                // 11'h3c7 :  DATA_OUT <= random_bits[30975:30944];
                // 11'h3c8 :  DATA_OUT <= random_bits[31007:30976];
                // 11'h3c9 :  DATA_OUT <= random_bits[31039:31008];
                // 11'h3ca :  DATA_OUT <= random_bits[31071:31040];
                // 11'h3cb :  DATA_OUT <= random_bits[31103:31072];
                // 11'h3cc :  DATA_OUT <= random_bits[31135:31104];
                // 11'h3cd :  DATA_OUT <= random_bits[31167:31136];
                // 11'h3ce :  DATA_OUT <= random_bits[31199:31168];
                // 11'h3cf :  DATA_OUT <= random_bits[31231:31200];
                // 11'h3d0 :  DATA_OUT <= random_bits[31263:31232];
                // 11'h3d1 :  DATA_OUT <= random_bits[31295:31264];
                // 11'h3d2 :  DATA_OUT <= random_bits[31327:31296];
                // 11'h3d3 :  DATA_OUT <= random_bits[31359:31328];
                // 11'h3d4 :  DATA_OUT <= random_bits[31391:31360];
                // 11'h3d5 :  DATA_OUT <= random_bits[31423:31392];
                // 11'h3d6 :  DATA_OUT <= random_bits[31455:31424];
                // 11'h3d7 :  DATA_OUT <= random_bits[31487:31456];
                // 11'h3d8 :  DATA_OUT <= random_bits[31519:31488];
                // 11'h3d9 :  DATA_OUT <= random_bits[31551:31520];
                // 11'h3da :  DATA_OUT <= random_bits[31583:31552];
                // 11'h3db :  DATA_OUT <= random_bits[31615:31584];
                // 11'h3dc :  DATA_OUT <= random_bits[31647:31616];
                // 11'h3dd :  DATA_OUT <= random_bits[31679:31648];
                // 11'h3de :  DATA_OUT <= random_bits[31711:31680];
                // 11'h3df :  DATA_OUT <= random_bits[31743:31712];
                // 11'h3e0 :  DATA_OUT <= random_bits[31775:31744];
                // 11'h3e1 :  DATA_OUT <= random_bits[31807:31776];
                // 11'h3e2 :  DATA_OUT <= random_bits[31839:31808];
                // 11'h3e3 :  DATA_OUT <= random_bits[31871:31840];
                // 11'h3e4 :  DATA_OUT <= random_bits[31903:31872];
                // 11'h3e5 :  DATA_OUT <= random_bits[31935:31904];
                // 11'h3e6 :  DATA_OUT <= random_bits[31967:31936];
                // 11'h3e7 :  DATA_OUT <= random_bits[31999:31968];
                // 11'h3e8 :  DATA_OUT <= random_bits[32031:32000];
                // 11'h3e9 :  DATA_OUT <= random_bits[32063:32032];
                // 11'h3ea :  DATA_OUT <= random_bits[32095:32064];
                // 11'h3eb :  DATA_OUT <= random_bits[32127:32096];
                // 11'h3ec :  DATA_OUT <= random_bits[32159:32128];
                // 11'h3ed :  DATA_OUT <= random_bits[32191:32160];
                // 11'h3ee :  DATA_OUT <= random_bits[32223:32192];
                // 11'h3ef :  DATA_OUT <= random_bits[32255:32224];
                // 11'h3f0 :  DATA_OUT <= random_bits[32287:32256];
                // 11'h3f1 :  DATA_OUT <= random_bits[32319:32288];
                // 11'h3f2 :  DATA_OUT <= random_bits[32351:32320];
                // 11'h3f3 :  DATA_OUT <= random_bits[32383:32352];
                // 11'h3f4 :  DATA_OUT <= random_bits[32415:32384];
                // 11'h3f5 :  DATA_OUT <= random_bits[32447:32416];
                // 11'h3f6 :  DATA_OUT <= random_bits[32479:32448];
                // 11'h3f7 :  DATA_OUT <= random_bits[32511:32480];
                // 11'h3f8 :  DATA_OUT <= random_bits[32543:32512];
                // 11'h3f9 :  DATA_OUT <= random_bits[32575:32544];
                // 11'h3fa :  DATA_OUT <= random_bits[32607:32576];
                // 11'h3fb :  DATA_OUT <= random_bits[32639:32608];
                // 11'h3fc :  DATA_OUT <= random_bits[32671:32640];
                // 11'h3fd :  DATA_OUT <= random_bits[32703:32672];
                // 11'h3fe :  DATA_OUT <= random_bits[32735:32704];
                // 11'h3ff :  DATA_OUT <= random_bits[32767:32736];
                
                //ZAPISYWANIE HASHA
                11'h400 :  DATA_OUT <= digest_data[31:0];
                11'h401 :  DATA_OUT <= digest_data[63:32];
                11'h402 :  DATA_OUT <= digest_data[91:64];
                11'h403 :  DATA_OUT <= digest_data[127:96];
                11'h404 :  DATA_OUT <= digest_data[159:128];
                11'h405 :  DATA_OUT <= digest_data[191:160];
                11'h406 :  DATA_OUT <= digest_data[223:192];
                11'h407 :  DATA_OUT <= digest_data[255:224];
                11'h408 :  DATA_OUT <= digest_data[287:256];
                11'h409 :  DATA_OUT <= digest_data[319:288];
                11'h40a :  DATA_OUT <= digest_data[351:320];
                11'h40b :  DATA_OUT <= digest_data[383:352];
                11'h40c :  DATA_OUT <= digest_data[415:384];
                11'h40d :  DATA_OUT <= digest_data[447:416];
                11'h40e :  DATA_OUT <= digest_data[479:448];
                11'h40f :  DATA_OUT <= digest_data[511:480];
                
                //ODCZYTAŁEM WSZYSTKO, PRZECHODZĘ W STAN reset
                11'h7ff :  state <= data_sended;
                
                default :  DATA_OUT <= random_bits[31:0];
            endcase
         end
         
         data_sended : begin
            ready <= 0;
            state <= reset;
         end
    endcase
    end
end
//assign sha3_din = random_bits[writed_words_counter*(32+1):writed_words_counter*32];

endmodule
